// Copyright 2009 Altera Corporation. All rights reserved.  
// Altera products are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.  
//
// This reference design file, and your use thereof, is subject to and governed
// by the terms and conditions of the applicable Altera Reference Design 
// License Agreement (either as signed by you or found at www.altera.com).  By
// using this reference design file, you indicate your acceptance of such terms
// and conditions between you and Altera Corporation.  In the event that you do
// not agree with such terms and conditions, you may not use the reference 
// design file and please promptly destroy any copies you have made.
//
// This reference design file is being provided on an "as-is" basis and as an 
// accommodation and therefore all warranties, representations or guarantees of 
// any kind (whether express, implied or statutory) including, without 
// limitation, warranties of merchantability, non-infringement, or fitness for
// a particular purpose, are specifically disclaimed.  By making this reference
// design file available, Altera expressly does not recommend, suggest or 
// require that this reference design file be used in combination with any 
// other product not provided by Altera.
/////////////////////////////////////////////////////////////////////////////

module font_rom (
    input clk,
    input [10:0] addr,
    output reg [23:0] out
);

reg [10:0] addr_r;
always @(posedge clk) begin
  addr_r <= addr;
  case (addr_r)
// rows 7 to 30
// start rec 0 h = 24 w = 22 ofs = 0
    11'd0 : out <= 24'b00001111111100000000000;
    11'd1 : out <= 24'b00001111111110000000000;
    11'd2 : out <= 24'b00001111111110000000000;
    11'd3 : out <= 24'b00000001111111000000000;
    11'd4 : out <= 24'b00000001111111000000000;
    11'd5 : out <= 24'b00000011110111100000000;
    11'd6 : out <= 24'b00000011110111100000000;
    11'd7 : out <= 24'b00000011100011100000000;
    11'd8 : out <= 24'b00000111100011110000000;
    11'd9 : out <= 24'b00000111000001110000000;
    11'd10 : out <= 24'b00001111000001111000000;
    11'd11 : out <= 24'b00001111111111111000000;
    11'd12 : out <= 24'b00011111111111111100000;
    11'd13 : out <= 24'b00011111111111111100000;
    11'd14 : out <= 24'b00111100000000011110000;
    11'd15 : out <= 24'b00111100000000011110000;
    11'd16 : out <= 24'b11111111000001111111100;
    11'd17 : out <= 24'b11111111000001111111100;
    11'd18 : out <= 24'b11111111000001111111100;
    11'd19 : out <= 24'b00000000000000000000000;
    11'd20 : out <= 24'b00000000000000000000000;
    11'd21 : out <= 24'b00000000000000000000000;
    11'd22 : out <= 24'b00000000000000000000000;
    11'd23 : out <= 24'b0;
    11'd24 : out <= 24'b0;
    11'd25 : out <= 24'b0;
    11'd26 : out <= 24'b0;

// start rec 1 h = 24 w = 19 ofs = 27
    11'd27 : out <= 24'b11111111111111000000000;
    11'd28 : out <= 24'b11111111111111110000000;
    11'd29 : out <= 24'b11111111111111110000000;
    11'd30 : out <= 24'b00011100000011111000000;
    11'd31 : out <= 24'b00011100000001111000000;
    11'd32 : out <= 24'b00011100000000111000000;
    11'd33 : out <= 24'b00011100000001111000000;
    11'd34 : out <= 24'b00011100000111111000000;
    11'd35 : out <= 24'b00011111111111110000000;
    11'd36 : out <= 24'b00011111111111110000000;
    11'd37 : out <= 24'b00011111111111111000000;
    11'd38 : out <= 24'b00011100000011111100000;
    11'd39 : out <= 24'b00011100000000111100000;
    11'd40 : out <= 24'b00011100000000111100000;
    11'd41 : out <= 24'b00011100000000011100000;
    11'd42 : out <= 24'b00011100000001111100000;
    11'd43 : out <= 24'b11111111111111111100000;
    11'd44 : out <= 24'b11111111111111111000000;
    11'd45 : out <= 24'b11111111111111110000000;
    11'd46 : out <= 24'b00000000000000000000000;
    11'd47 : out <= 24'b00000000000000000000000;
    11'd48 : out <= 24'b00000000000000000000000;
    11'd49 : out <= 24'b00000000000000000000000;
    11'd50 : out <= 24'b0;
    11'd51 : out <= 24'b0;
    11'd52 : out <= 24'b0;
    11'd53 : out <= 24'b0;

// start rec 2 h = 24 w = 18 ofs = 54
    11'd54 : out <= 24'b00000111111111111000000;
    11'd55 : out <= 24'b00011111111111111000000;
    11'd56 : out <= 24'b00111111111111111000000;
    11'd57 : out <= 24'b01111111001111111000000;
    11'd58 : out <= 24'b01111100000001111000000;
    11'd59 : out <= 24'b11111000000000111000000;
    11'd60 : out <= 24'b11110000000000111000000;
    11'd61 : out <= 24'b11110000000000000000000;
    11'd62 : out <= 24'b11100000000000000000000;
    11'd63 : out <= 24'b11100000000000000000000;
    11'd64 : out <= 24'b11100000000000000000000;
    11'd65 : out <= 24'b11100000000000000000000;
    11'd66 : out <= 24'b11110000000000000000000;
    11'd67 : out <= 24'b11110000000000111000000;
    11'd68 : out <= 24'b01111000000001111000000;
    11'd69 : out <= 24'b01111111000111111000000;
    11'd70 : out <= 24'b00111111111111111000000;
    11'd71 : out <= 24'b00011111111111110000000;
    11'd72 : out <= 24'b00000111111111000000000;
    11'd73 : out <= 24'b00000000000000000000000;
    11'd74 : out <= 24'b00000000000000000000000;
    11'd75 : out <= 24'b00000000000000000000000;
    11'd76 : out <= 24'b00000000000000000000000;
    11'd77 : out <= 24'b0;
    11'd78 : out <= 24'b0;
    11'd79 : out <= 24'b0;
    11'd80 : out <= 24'b0;

// start rec 3 h = 24 w = 18 ofs = 81
    11'd81 : out <= 24'b11111111111100000000000;
    11'd82 : out <= 24'b11111111111111000000000;
    11'd83 : out <= 24'b11111111111111100000000;
    11'd84 : out <= 24'b00111000001111110000000;
    11'd85 : out <= 24'b00111000000011110000000;
    11'd86 : out <= 24'b00111000000001111000000;
    11'd87 : out <= 24'b00111000000001111000000;
    11'd88 : out <= 24'b00111000000001111000000;
    11'd89 : out <= 24'b00111000000000111000000;
    11'd90 : out <= 24'b00111000000000111000000;
    11'd91 : out <= 24'b00111000000000111000000;
    11'd92 : out <= 24'b00111000000000111000000;
    11'd93 : out <= 24'b00111000000001111000000;
    11'd94 : out <= 24'b00111000000001111000000;
    11'd95 : out <= 24'b00111000000011111000000;
    11'd96 : out <= 24'b00111000001111110000000;
    11'd97 : out <= 24'b11111111111111100000000;
    11'd98 : out <= 24'b11111111111111000000000;
    11'd99 : out <= 24'b11111111111110000000000;
    11'd100 : out <= 24'b00000000000000000000000;
    11'd101 : out <= 24'b00000000000000000000000;
    11'd102 : out <= 24'b00000000000000000000000;
    11'd103 : out <= 24'b00000000000000000000000;
    11'd104 : out <= 24'b0;
    11'd105 : out <= 24'b0;
    11'd106 : out <= 24'b0;
    11'd107 : out <= 24'b0;

// start rec 4 h = 24 w = 18 ofs = 108
    11'd108 : out <= 24'b11111111111111110000000;
    11'd109 : out <= 24'b11111111111111110000000;
    11'd110 : out <= 24'b11111111111111110000000;
    11'd111 : out <= 24'b00011100000001110000000;
    11'd112 : out <= 24'b00011100000001110000000;
    11'd113 : out <= 24'b00011100000001110000000;
    11'd114 : out <= 24'b00011100011101110000000;
    11'd115 : out <= 24'b00011100011100000000000;
    11'd116 : out <= 24'b00011111111100000000000;
    11'd117 : out <= 24'b00011111111100000000000;
    11'd118 : out <= 24'b00011111111100000000000;
    11'd119 : out <= 24'b00011100011100000000000;
    11'd120 : out <= 24'b00011100011100111000000;
    11'd121 : out <= 24'b00011100000000111000000;
    11'd122 : out <= 24'b00011100000000111000000;
    11'd123 : out <= 24'b00011100000000111000000;
    11'd124 : out <= 24'b11111111111111111000000;
    11'd125 : out <= 24'b11111111111111111000000;
    11'd126 : out <= 24'b11111111111111111000000;
    11'd127 : out <= 24'b00000000000000000000000;
    11'd128 : out <= 24'b00000000000000000000000;
    11'd129 : out <= 24'b00000000000000000000000;
    11'd130 : out <= 24'b00000000000000000000000;
    11'd131 : out <= 24'b0;
    11'd132 : out <= 24'b0;
    11'd133 : out <= 24'b0;
    11'd134 : out <= 24'b0;

// start rec 5 h = 24 w = 18 ofs = 135
    11'd135 : out <= 24'b11111111111111111000000;
    11'd136 : out <= 24'b11111111111111111000000;
    11'd137 : out <= 24'b11111111111111111000000;
    11'd138 : out <= 24'b00011100000000111000000;
    11'd139 : out <= 24'b00011100000000111000000;
    11'd140 : out <= 24'b00011100000000111000000;
    11'd141 : out <= 24'b00011100011100111000000;
    11'd142 : out <= 24'b00011100011100000000000;
    11'd143 : out <= 24'b00011111111100000000000;
    11'd144 : out <= 24'b00011111111100000000000;
    11'd145 : out <= 24'b00011111111100000000000;
    11'd146 : out <= 24'b00011100011100000000000;
    11'd147 : out <= 24'b00011100011100000000000;
    11'd148 : out <= 24'b00011100000000000000000;
    11'd149 : out <= 24'b00011100000000000000000;
    11'd150 : out <= 24'b00011100000000000000000;
    11'd151 : out <= 24'b11111111111000000000000;
    11'd152 : out <= 24'b11111111111000000000000;
    11'd153 : out <= 24'b11111111111000000000000;
    11'd154 : out <= 24'b00000000000000000000000;
    11'd155 : out <= 24'b00000000000000000000000;
    11'd156 : out <= 24'b00000000000000000000000;
    11'd157 : out <= 24'b00000000000000000000000;
    11'd158 : out <= 24'b0;
    11'd159 : out <= 24'b0;
    11'd160 : out <= 24'b0;
    11'd161 : out <= 24'b0;

// start rec 6 h = 24 w = 19 ofs = 162
    11'd162 : out <= 24'b00001111111111110000000;
    11'd163 : out <= 24'b00011111111111110000000;
    11'd164 : out <= 24'b00111111111111110000000;
    11'd165 : out <= 24'b01111110001111110000000;
    11'd166 : out <= 24'b01111000000011110000000;
    11'd167 : out <= 24'b11110000000011110000000;
    11'd168 : out <= 24'b11110000000000000000000;
    11'd169 : out <= 24'b11110000000000000000000;
    11'd170 : out <= 24'b11100000000000000000000;
    11'd171 : out <= 24'b11100000111111111100000;
    11'd172 : out <= 24'b11100000111111111100000;
    11'd173 : out <= 24'b11100000111111111100000;
    11'd174 : out <= 24'b11110000000001110000000;
    11'd175 : out <= 24'b11110000000001110000000;
    11'd176 : out <= 24'b11111000000011110000000;
    11'd177 : out <= 24'b01111110001111110000000;
    11'd178 : out <= 24'b00111111111111110000000;
    11'd179 : out <= 24'b00011111111111100000000;
    11'd180 : out <= 24'b00001111111110000000000;
    11'd181 : out <= 24'b00000000000000000000000;
    11'd182 : out <= 24'b00000000000000000000000;
    11'd183 : out <= 24'b00000000000000000000000;
    11'd184 : out <= 24'b00000000000000000000000;
    11'd185 : out <= 24'b0;
    11'd186 : out <= 24'b0;
    11'd187 : out <= 24'b0;
    11'd188 : out <= 24'b0;

// start rec 7 h = 24 w = 18 ofs = 189
    11'd189 : out <= 24'b11111110001111111000000;
    11'd190 : out <= 24'b11111110001111111000000;
    11'd191 : out <= 24'b11111110001111111000000;
    11'd192 : out <= 24'b00111000000011100000000;
    11'd193 : out <= 24'b00111000000011100000000;
    11'd194 : out <= 24'b00111000000011100000000;
    11'd195 : out <= 24'b00111000000011100000000;
    11'd196 : out <= 24'b00111000000011100000000;
    11'd197 : out <= 24'b00111111111111100000000;
    11'd198 : out <= 24'b00111111111111100000000;
    11'd199 : out <= 24'b00111111111111100000000;
    11'd200 : out <= 24'b00111000000011100000000;
    11'd201 : out <= 24'b00111000000011100000000;
    11'd202 : out <= 24'b00111000000011100000000;
    11'd203 : out <= 24'b00111000000011100000000;
    11'd204 : out <= 24'b00111000000011100000000;
    11'd205 : out <= 24'b11111110001111111000000;
    11'd206 : out <= 24'b11111110001111111000000;
    11'd207 : out <= 24'b11111110001111111000000;
    11'd208 : out <= 24'b00000000000000000000000;
    11'd209 : out <= 24'b00000000000000000000000;
    11'd210 : out <= 24'b00000000000000000000000;
    11'd211 : out <= 24'b00000000000000000000000;
    11'd212 : out <= 24'b0;
    11'd213 : out <= 24'b0;
    11'd214 : out <= 24'b0;
    11'd215 : out <= 24'b0;

// start rec 8 h = 24 w = 14 ofs = 216
    11'd216 : out <= 24'b11111111111110000000000;
    11'd217 : out <= 24'b11111111111110000000000;
    11'd218 : out <= 24'b11111111111110000000000;
    11'd219 : out <= 24'b00000111000000000000000;
    11'd220 : out <= 24'b00000111000000000000000;
    11'd221 : out <= 24'b00000111000000000000000;
    11'd222 : out <= 24'b00000111000000000000000;
    11'd223 : out <= 24'b00000111000000000000000;
    11'd224 : out <= 24'b00000111000000000000000;
    11'd225 : out <= 24'b00000111000000000000000;
    11'd226 : out <= 24'b00000111000000000000000;
    11'd227 : out <= 24'b00000111000000000000000;
    11'd228 : out <= 24'b00000111000000000000000;
    11'd229 : out <= 24'b00000111000000000000000;
    11'd230 : out <= 24'b00000111000000000000000;
    11'd231 : out <= 24'b00000111000000000000000;
    11'd232 : out <= 24'b11111111111110000000000;
    11'd233 : out <= 24'b11111111111110000000000;
    11'd234 : out <= 24'b11111111111110000000000;
    11'd235 : out <= 24'b00000000000000000000000;
    11'd236 : out <= 24'b00000000000000000000000;
    11'd237 : out <= 24'b00000000000000000000000;
    11'd238 : out <= 24'b00000000000000000000000;
    11'd239 : out <= 24'b0;
    11'd240 : out <= 24'b0;
    11'd241 : out <= 24'b0;
    11'd242 : out <= 24'b0;

// start rec 9 h = 24 w = 18 ofs = 243
    11'd243 : out <= 24'b00001111111111111000000;
    11'd244 : out <= 24'b00001111111111111000000;
    11'd245 : out <= 24'b00001111111111111000000;
    11'd246 : out <= 24'b00000000001110000000000;
    11'd247 : out <= 24'b00000000001110000000000;
    11'd248 : out <= 24'b00000000001110000000000;
    11'd249 : out <= 24'b00000000001110000000000;
    11'd250 : out <= 24'b00000000001110000000000;
    11'd251 : out <= 24'b00000000001110000000000;
    11'd252 : out <= 24'b00000000001110000000000;
    11'd253 : out <= 24'b11100000001110000000000;
    11'd254 : out <= 24'b11100000001110000000000;
    11'd255 : out <= 24'b11100000001110000000000;
    11'd256 : out <= 24'b11100000001110000000000;
    11'd257 : out <= 24'b11100000011110000000000;
    11'd258 : out <= 24'b11111101111110000000000;
    11'd259 : out <= 24'b11111111111100000000000;
    11'd260 : out <= 24'b11111111111000000000000;
    11'd261 : out <= 24'b00111111110000000000000;
    11'd262 : out <= 24'b00000000000000000000000;
    11'd263 : out <= 24'b00000000000000000000000;
    11'd264 : out <= 24'b00000000000000000000000;
    11'd265 : out <= 24'b00000000000000000000000;
    11'd266 : out <= 24'b0;
    11'd267 : out <= 24'b0;
    11'd268 : out <= 24'b0;
    11'd269 : out <= 24'b0;

// start rec 10 h = 24 w = 20 ofs = 270
    11'd270 : out <= 24'b11111111100011111110000;
    11'd271 : out <= 24'b11111111100011111110000;
    11'd272 : out <= 24'b11111111100011111110000;
    11'd273 : out <= 24'b00011100000111110000000;
    11'd274 : out <= 24'b00011100001111100000000;
    11'd275 : out <= 24'b00011100011111000000000;
    11'd276 : out <= 24'b00011101111100000000000;
    11'd277 : out <= 24'b00011111111000000000000;
    11'd278 : out <= 24'b00011111111100000000000;
    11'd279 : out <= 24'b00011111111110000000000;
    11'd280 : out <= 24'b00011110011111000000000;
    11'd281 : out <= 24'b00011100001111000000000;
    11'd282 : out <= 24'b00011100000111100000000;
    11'd283 : out <= 24'b00011100000111100000000;
    11'd284 : out <= 24'b00011100000011110000000;
    11'd285 : out <= 24'b00011100000011110000000;
    11'd286 : out <= 24'b11111111100001111110000;
    11'd287 : out <= 24'b11111111100001111110000;
    11'd288 : out <= 24'b11111111100001111110000;
    11'd289 : out <= 24'b00000000000000000000000;
    11'd290 : out <= 24'b00000000000000000000000;
    11'd291 : out <= 24'b00000000000000000000000;
    11'd292 : out <= 24'b00000000000000000000000;
    11'd293 : out <= 24'b0;
    11'd294 : out <= 24'b0;
    11'd295 : out <= 24'b0;
    11'd296 : out <= 24'b0;

// start rec 11 h = 24 w = 18 ofs = 297
    11'd297 : out <= 24'b11111111111000000000000;
    11'd298 : out <= 24'b11111111111000000000000;
    11'd299 : out <= 24'b11111111111000000000000;
    11'd300 : out <= 24'b00001110000000000000000;
    11'd301 : out <= 24'b00001110000000000000000;
    11'd302 : out <= 24'b00001110000000000000000;
    11'd303 : out <= 24'b00001110000000000000000;
    11'd304 : out <= 24'b00001110000000000000000;
    11'd305 : out <= 24'b00001110000000000000000;
    11'd306 : out <= 24'b00001110000000000000000;
    11'd307 : out <= 24'b00001110000000000000000;
    11'd308 : out <= 24'b00001110000000111000000;
    11'd309 : out <= 24'b00001110000000111000000;
    11'd310 : out <= 24'b00001110000000111000000;
    11'd311 : out <= 24'b00001110000000111000000;
    11'd312 : out <= 24'b00001110000000111000000;
    11'd313 : out <= 24'b11111111111111111000000;
    11'd314 : out <= 24'b11111111111111111000000;
    11'd315 : out <= 24'b11111111111111111000000;
    11'd316 : out <= 24'b00000000000000000000000;
    11'd317 : out <= 24'b00000000000000000000000;
    11'd318 : out <= 24'b00000000000000000000000;
    11'd319 : out <= 24'b00000000000000000000000;
    11'd320 : out <= 24'b0;
    11'd321 : out <= 24'b0;
    11'd322 : out <= 24'b0;
    11'd323 : out <= 24'b0;

// start rec 12 h = 24 w = 22 ofs = 324
    11'd324 : out <= 24'b11111100000000011111100;
    11'd325 : out <= 24'b11111100000000011111100;
    11'd326 : out <= 24'b11111110000000111111100;
    11'd327 : out <= 24'b00111110000000111110000;
    11'd328 : out <= 24'b00111111000001111110000;
    11'd329 : out <= 24'b00111111000001111110000;
    11'd330 : out <= 24'b00111111100011111110000;
    11'd331 : out <= 24'b00111011110111101110000;
    11'd332 : out <= 24'b00111011110111101110000;
    11'd333 : out <= 24'b00111001111111001110000;
    11'd334 : out <= 24'b00111001111111001110000;
    11'd335 : out <= 24'b00111000111110001110000;
    11'd336 : out <= 24'b00111000111110001110000;
    11'd337 : out <= 24'b00111000011100001110000;
    11'd338 : out <= 24'b00111000011100001110000;
    11'd339 : out <= 24'b00111000000000001110000;
    11'd340 : out <= 24'b11111111000001111111100;
    11'd341 : out <= 24'b11111111000001111111100;
    11'd342 : out <= 24'b11111111000001111111100;
    11'd343 : out <= 24'b00000000000000000000000;
    11'd344 : out <= 24'b00000000000000000000000;
    11'd345 : out <= 24'b00000000000000000000000;
    11'd346 : out <= 24'b00000000000000000000000;
    11'd347 : out <= 24'b0;
    11'd348 : out <= 24'b0;
    11'd349 : out <= 24'b0;
    11'd350 : out <= 24'b0;

// start rec 13 h = 24 w = 20 ofs = 351
    11'd351 : out <= 24'b11111100000111111110000;
    11'd352 : out <= 24'b11111110000111111110000;
    11'd353 : out <= 24'b11111110000111111110000;
    11'd354 : out <= 24'b00011111000000111000000;
    11'd355 : out <= 24'b00011111100000111000000;
    11'd356 : out <= 24'b00011111100000111000000;
    11'd357 : out <= 24'b00011111110000111000000;
    11'd358 : out <= 24'b00011101111000111000000;
    11'd359 : out <= 24'b00011101111000111000000;
    11'd360 : out <= 24'b00011100111100111000000;
    11'd361 : out <= 24'b00011100011110111000000;
    11'd362 : out <= 24'b00011100011111111000000;
    11'd363 : out <= 24'b00011100001111111000000;
    11'd364 : out <= 24'b00011100000111111000000;
    11'd365 : out <= 24'b00011100000111111000000;
    11'd366 : out <= 24'b00011100000011111000000;
    11'd367 : out <= 24'b01111111100001111000000;
    11'd368 : out <= 24'b01111111100001111000000;
    11'd369 : out <= 24'b01111111100000111000000;
    11'd370 : out <= 24'b00000000000000000000000;
    11'd371 : out <= 24'b00000000000000000000000;
    11'd372 : out <= 24'b00000000000000000000000;
    11'd373 : out <= 24'b00000000000000000000000;
    11'd374 : out <= 24'b0;
    11'd375 : out <= 24'b0;
    11'd376 : out <= 24'b0;
    11'd377 : out <= 24'b0;

// start rec 14 h = 24 w = 18 ofs = 378
    11'd378 : out <= 24'b00000111111100000000000;
    11'd379 : out <= 24'b00011111111111000000000;
    11'd380 : out <= 24'b00111111111111100000000;
    11'd381 : out <= 24'b01111111011111110000000;
    11'd382 : out <= 24'b01111100000111110000000;
    11'd383 : out <= 24'b11111000000011111000000;
    11'd384 : out <= 24'b11110000000001111000000;
    11'd385 : out <= 24'b11110000000001111000000;
    11'd386 : out <= 24'b11100000000000111000000;
    11'd387 : out <= 24'b11100000000000111000000;
    11'd388 : out <= 24'b11100000000000111000000;
    11'd389 : out <= 24'b11110000000001111000000;
    11'd390 : out <= 24'b11110000000001111000000;
    11'd391 : out <= 24'b11111000000011111000000;
    11'd392 : out <= 24'b01111100000111110000000;
    11'd393 : out <= 24'b01111111011111110000000;
    11'd394 : out <= 24'b00111111111111100000000;
    11'd395 : out <= 24'b00011111111111000000000;
    11'd396 : out <= 24'b00000111111100000000000;
    11'd397 : out <= 24'b00000000000000000000000;
    11'd398 : out <= 24'b00000000000000000000000;
    11'd399 : out <= 24'b00000000000000000000000;
    11'd400 : out <= 24'b00000000000000000000000;
    11'd401 : out <= 24'b0;
    11'd402 : out <= 24'b0;
    11'd403 : out <= 24'b0;
    11'd404 : out <= 24'b0;

// start rec 15 h = 24 w = 18 ofs = 405
    11'd405 : out <= 24'b11111111111111000000000;
    11'd406 : out <= 24'b11111111111111100000000;
    11'd407 : out <= 24'b11111111111111110000000;
    11'd408 : out <= 24'b00011100000111111000000;
    11'd409 : out <= 24'b00011100000001111000000;
    11'd410 : out <= 24'b00011100000001111000000;
    11'd411 : out <= 24'b00011100000000111000000;
    11'd412 : out <= 24'b00011100000001111000000;
    11'd413 : out <= 24'b00011100000001111000000;
    11'd414 : out <= 24'b00011100001111111000000;
    11'd415 : out <= 24'b00011111111111110000000;
    11'd416 : out <= 24'b00011111111111100000000;
    11'd417 : out <= 24'b00011111111110000000000;
    11'd418 : out <= 24'b00011100000000000000000;
    11'd419 : out <= 24'b00011100000000000000000;
    11'd420 : out <= 24'b00011100000000000000000;
    11'd421 : out <= 24'b11111111111000000000000;
    11'd422 : out <= 24'b11111111111000000000000;
    11'd423 : out <= 24'b11111111111000000000000;
    11'd424 : out <= 24'b00000000000000000000000;
    11'd425 : out <= 24'b00000000000000000000000;
    11'd426 : out <= 24'b00000000000000000000000;
    11'd427 : out <= 24'b00000000000000000000000;
    11'd428 : out <= 24'b0;
    11'd429 : out <= 24'b0;
    11'd430 : out <= 24'b0;
    11'd431 : out <= 24'b0;

// start rec 16 h = 24 w = 18 ofs = 432
    11'd432 : out <= 24'b00000111111100000000000;
    11'd433 : out <= 24'b00011111111111000000000;
    11'd434 : out <= 24'b00111111111111100000000;
    11'd435 : out <= 24'b00111111011111110000000;
    11'd436 : out <= 24'b01111100000111110000000;
    11'd437 : out <= 24'b11111000000011111000000;
    11'd438 : out <= 24'b11110000000001111000000;
    11'd439 : out <= 24'b11110000000001111000000;
    11'd440 : out <= 24'b11100000000000111000000;
    11'd441 : out <= 24'b11100000000000111000000;
    11'd442 : out <= 24'b11100000000000111000000;
    11'd443 : out <= 24'b11110000000001111000000;
    11'd444 : out <= 24'b11110000000001111000000;
    11'd445 : out <= 24'b11111000000011111000000;
    11'd446 : out <= 24'b01111100000111110000000;
    11'd447 : out <= 24'b01111111011111110000000;
    11'd448 : out <= 24'b00111111111111100000000;
    11'd449 : out <= 24'b00011111111111000000000;
    11'd450 : out <= 24'b00001111111100000000000;
    11'd451 : out <= 24'b00000111111111111000000;
    11'd452 : out <= 24'b00011111111111111000000;
    11'd453 : out <= 24'b00011111111111111000000;
    11'd454 : out <= 24'b00011111001111110000000;
    11'd455 : out <= 24'b0;
    11'd456 : out <= 24'b0;
    11'd457 : out <= 24'b0;
    11'd458 : out <= 24'b0;

// start rec 17 h = 24 w = 21 ofs = 459
    11'd459 : out <= 24'b11111111111111000000000;
    11'd460 : out <= 24'b11111111111111100000000;
    11'd461 : out <= 24'b11111111111111110000000;
    11'd462 : out <= 24'b00011100000111111000000;
    11'd463 : out <= 24'b00011100000001111000000;
    11'd464 : out <= 24'b00011100000000111000000;
    11'd465 : out <= 24'b00011100000001111000000;
    11'd466 : out <= 24'b00011100000001111000000;
    11'd467 : out <= 24'b00011100001111111000000;
    11'd468 : out <= 24'b00011111111111110000000;
    11'd469 : out <= 24'b00011111111111100000000;
    11'd470 : out <= 24'b00011111111111100000000;
    11'd471 : out <= 24'b00011100001111110000000;
    11'd472 : out <= 24'b00011100000111111000000;
    11'd473 : out <= 24'b00011100000011111000000;
    11'd474 : out <= 24'b00011100000001111100000;
    11'd475 : out <= 24'b11111111100000111111000;
    11'd476 : out <= 24'b11111111100000011111000;
    11'd477 : out <= 24'b11111111100000011111000;
    11'd478 : out <= 24'b00000000000000000000000;
    11'd479 : out <= 24'b00000000000000000000000;
    11'd480 : out <= 24'b00000000000000000000000;
    11'd481 : out <= 24'b00000000000000000000000;
    11'd482 : out <= 24'b0;
    11'd483 : out <= 24'b0;
    11'd484 : out <= 24'b0;
    11'd485 : out <= 24'b0;

// start rec 18 h = 24 w = 16 ofs = 486
    11'd486 : out <= 24'b00001111111111000000000;
    11'd487 : out <= 24'b00111111111111000000000;
    11'd488 : out <= 24'b00111111111111000000000;
    11'd489 : out <= 24'b01111110011111000000000;
    11'd490 : out <= 24'b01111000000111000000000;
    11'd491 : out <= 24'b01110000000111000000000;
    11'd492 : out <= 24'b01111000000111000000000;
    11'd493 : out <= 24'b01111111000000000000000;
    11'd494 : out <= 24'b00111111111100000000000;
    11'd495 : out <= 24'b00111111111111000000000;
    11'd496 : out <= 24'b00001111111111000000000;
    11'd497 : out <= 24'b00000000111111100000000;
    11'd498 : out <= 24'b00000000000111100000000;
    11'd499 : out <= 24'b11100000000011100000000;
    11'd500 : out <= 24'b11100000000111100000000;
    11'd501 : out <= 24'b11111100011111100000000;
    11'd502 : out <= 24'b11111111111111100000000;
    11'd503 : out <= 24'b11111111111111000000000;
    11'd504 : out <= 24'b11111111111100000000000;
    11'd505 : out <= 24'b00000000000000000000000;
    11'd506 : out <= 24'b00000000000000000000000;
    11'd507 : out <= 24'b00000000000000000000000;
    11'd508 : out <= 24'b00000000000000000000000;
    11'd509 : out <= 24'b0;
    11'd510 : out <= 24'b0;
    11'd511 : out <= 24'b0;
    11'd512 : out <= 24'b0;

// start rec 19 h = 24 w = 18 ofs = 513
    11'd513 : out <= 24'b11111111111111111000000;
    11'd514 : out <= 24'b11111111111111111000000;
    11'd515 : out <= 24'b11111111111111111000000;
    11'd516 : out <= 24'b11100001110000111000000;
    11'd517 : out <= 24'b11100001110000111000000;
    11'd518 : out <= 24'b11100001110000111000000;
    11'd519 : out <= 24'b11100001110000111000000;
    11'd520 : out <= 24'b11100001110000111000000;
    11'd521 : out <= 24'b00000001110000000000000;
    11'd522 : out <= 24'b00000001110000000000000;
    11'd523 : out <= 24'b00000001110000000000000;
    11'd524 : out <= 24'b00000001110000000000000;
    11'd525 : out <= 24'b00000001110000000000000;
    11'd526 : out <= 24'b00000001110000000000000;
    11'd527 : out <= 24'b00000001110000000000000;
    11'd528 : out <= 24'b00000001110000000000000;
    11'd529 : out <= 24'b00011111111111000000000;
    11'd530 : out <= 24'b00011111111111000000000;
    11'd531 : out <= 24'b00011111111111000000000;
    11'd532 : out <= 24'b00000000000000000000000;
    11'd533 : out <= 24'b00000000000000000000000;
    11'd534 : out <= 24'b00000000000000000000000;
    11'd535 : out <= 24'b00000000000000000000000;
    11'd536 : out <= 24'b0;
    11'd537 : out <= 24'b0;
    11'd538 : out <= 24'b0;
    11'd539 : out <= 24'b0;

// start rec 20 h = 24 w = 20 ofs = 540
    11'd540 : out <= 24'b11111111000111111110000;
    11'd541 : out <= 24'b11111111000111111110000;
    11'd542 : out <= 24'b11111111000111111110000;
    11'd543 : out <= 24'b00111000000000111000000;
    11'd544 : out <= 24'b00111000000000111000000;
    11'd545 : out <= 24'b00111000000000111000000;
    11'd546 : out <= 24'b00111000000000111000000;
    11'd547 : out <= 24'b00111000000000111000000;
    11'd548 : out <= 24'b00111000000000111000000;
    11'd549 : out <= 24'b00111000000000111000000;
    11'd550 : out <= 24'b00111000000000111000000;
    11'd551 : out <= 24'b00111000000000111000000;
    11'd552 : out <= 24'b00111000000000111000000;
    11'd553 : out <= 24'b00111100000001111000000;
    11'd554 : out <= 24'b00111100000001111000000;
    11'd555 : out <= 24'b00011111000111110000000;
    11'd556 : out <= 24'b00011111111111110000000;
    11'd557 : out <= 24'b00001111111111100000000;
    11'd558 : out <= 24'b00000011111110000000000;
    11'd559 : out <= 24'b00000000000000000000000;
    11'd560 : out <= 24'b00000000000000000000000;
    11'd561 : out <= 24'b00000000000000000000000;
    11'd562 : out <= 24'b00000000000000000000000;
    11'd563 : out <= 24'b0;
    11'd564 : out <= 24'b0;
    11'd565 : out <= 24'b0;
    11'd566 : out <= 24'b0;

// start rec 21 h = 24 w = 22 ofs = 567
    11'd567 : out <= 24'b11111111000001111111100;
    11'd568 : out <= 24'b11111111000001111111100;
    11'd569 : out <= 24'b11111111000001111111100;
    11'd570 : out <= 24'b00111100000000011110000;
    11'd571 : out <= 24'b00111100000000011110000;
    11'd572 : out <= 24'b00011110000000111100000;
    11'd573 : out <= 24'b00011110000000111100000;
    11'd574 : out <= 24'b00001111000001111000000;
    11'd575 : out <= 24'b00001111000001111000000;
    11'd576 : out <= 24'b00000111100011110000000;
    11'd577 : out <= 24'b00000111100011110000000;
    11'd578 : out <= 24'b00000111110111100000000;
    11'd579 : out <= 24'b00000011110111100000000;
    11'd580 : out <= 24'b00000011111111100000000;
    11'd581 : out <= 24'b00000001111111000000000;
    11'd582 : out <= 24'b00000001111111000000000;
    11'd583 : out <= 24'b00000000111110000000000;
    11'd584 : out <= 24'b00000000111110000000000;
    11'd585 : out <= 24'b00000000011100000000000;
    11'd586 : out <= 24'b00000000000000000000000;
    11'd587 : out <= 24'b00000000000000000000000;
    11'd588 : out <= 24'b00000000000000000000000;
    11'd589 : out <= 24'b00000000000000000000000;
    11'd590 : out <= 24'b0;
    11'd591 : out <= 24'b0;
    11'd592 : out <= 24'b0;
    11'd593 : out <= 24'b0;

// start rec 22 h = 24 w = 22 ofs = 594
    11'd594 : out <= 24'b11111111100011111111100;
    11'd595 : out <= 24'b11111111100011111111100;
    11'd596 : out <= 24'b11111111100011111111100;
    11'd597 : out <= 24'b00111100000000011110000;
    11'd598 : out <= 24'b00111100000000011110000;
    11'd599 : out <= 24'b00111100011100011110000;
    11'd600 : out <= 24'b00111100011100011110000;
    11'd601 : out <= 24'b00111100111110011110000;
    11'd602 : out <= 24'b00111100111110011110000;
    11'd603 : out <= 24'b00011100111110011100000;
    11'd604 : out <= 24'b00011111110111111100000;
    11'd605 : out <= 24'b00011111110111111100000;
    11'd606 : out <= 24'b00011111110111111100000;
    11'd607 : out <= 24'b00011111100011111100000;
    11'd608 : out <= 24'b00011111100011111100000;
    11'd609 : out <= 24'b00011111100011111100000;
    11'd610 : out <= 24'b00001111000001111000000;
    11'd611 : out <= 24'b00001111000001111000000;
    11'd612 : out <= 24'b00001110000000111000000;
    11'd613 : out <= 24'b00000000000000000000000;
    11'd614 : out <= 24'b00000000000000000000000;
    11'd615 : out <= 24'b00000000000000000000000;
    11'd616 : out <= 24'b00000000000000000000000;
    11'd617 : out <= 24'b0;
    11'd618 : out <= 24'b0;
    11'd619 : out <= 24'b0;
    11'd620 : out <= 24'b0;

// start rec 23 h = 24 w = 20 ofs = 621
    11'd621 : out <= 24'b11111110000011111110000;
    11'd622 : out <= 24'b11111110000011111110000;
    11'd623 : out <= 24'b11111110000011111110000;
    11'd624 : out <= 24'b00111100000001111000000;
    11'd625 : out <= 24'b00011110000011110000000;
    11'd626 : out <= 24'b00001111000111100000000;
    11'd627 : out <= 24'b00000111101111000000000;
    11'd628 : out <= 24'b00000011111110000000000;
    11'd629 : out <= 24'b00000001111100000000000;
    11'd630 : out <= 24'b00000001111100000000000;
    11'd631 : out <= 24'b00000001111100000000000;
    11'd632 : out <= 24'b00000011111110000000000;
    11'd633 : out <= 24'b00000111101111000000000;
    11'd634 : out <= 24'b00001111000111100000000;
    11'd635 : out <= 24'b00011110000011110000000;
    11'd636 : out <= 24'b00111100000001111000000;
    11'd637 : out <= 24'b11111110000011111110000;
    11'd638 : out <= 24'b11111110000011111110000;
    11'd639 : out <= 24'b11111110000011111110000;
    11'd640 : out <= 24'b00000000000000000000000;
    11'd641 : out <= 24'b00000000000000000000000;
    11'd642 : out <= 24'b00000000000000000000000;
    11'd643 : out <= 24'b00000000000000000000000;
    11'd644 : out <= 24'b0;
    11'd645 : out <= 24'b0;
    11'd646 : out <= 24'b0;
    11'd647 : out <= 24'b0;

// start rec 24 h = 24 w = 18 ofs = 648
    11'd648 : out <= 24'b11111110001111111000000;
    11'd649 : out <= 24'b11111110001111111000000;
    11'd650 : out <= 24'b11111110001111111000000;
    11'd651 : out <= 24'b00111100000111100000000;
    11'd652 : out <= 24'b00111100000111100000000;
    11'd653 : out <= 24'b00011110001111000000000;
    11'd654 : out <= 24'b00001111011110000000000;
    11'd655 : out <= 24'b00001111011110000000000;
    11'd656 : out <= 24'b00000111111100000000000;
    11'd657 : out <= 24'b00000011111000000000000;
    11'd658 : out <= 24'b00000011111000000000000;
    11'd659 : out <= 24'b00000001110000000000000;
    11'd660 : out <= 24'b00000001110000000000000;
    11'd661 : out <= 24'b00000001110000000000000;
    11'd662 : out <= 24'b00000001110000000000000;
    11'd663 : out <= 24'b00000001110000000000000;
    11'd664 : out <= 24'b00011111111111000000000;
    11'd665 : out <= 24'b00011111111111000000000;
    11'd666 : out <= 24'b00011111111111000000000;
    11'd667 : out <= 24'b00000000000000000000000;
    11'd668 : out <= 24'b00000000000000000000000;
    11'd669 : out <= 24'b00000000000000000000000;
    11'd670 : out <= 24'b00000000000000000000000;
    11'd671 : out <= 24'b0;
    11'd672 : out <= 24'b0;
    11'd673 : out <= 24'b0;
    11'd674 : out <= 24'b0;

// start rec 25 h = 24 w = 16 ofs = 675
    11'd675 : out <= 24'b01111111111111000000000;
    11'd676 : out <= 24'b01111111111111000000000;
    11'd677 : out <= 24'b01111111111111000000000;
    11'd678 : out <= 24'b01110000001111000000000;
    11'd679 : out <= 24'b01110000011110000000000;
    11'd680 : out <= 24'b01110000111100000000000;
    11'd681 : out <= 24'b01110000111100000000000;
    11'd682 : out <= 24'b00000001111000000000000;
    11'd683 : out <= 24'b00000011110000000000000;
    11'd684 : out <= 24'b00000111100000000000000;
    11'd685 : out <= 24'b00001111000000000000000;
    11'd686 : out <= 24'b00011110000000000000000;
    11'd687 : out <= 24'b00111100000011100000000;
    11'd688 : out <= 24'b00111100000011100000000;
    11'd689 : out <= 24'b01111000000011100000000;
    11'd690 : out <= 24'b11110000000011100000000;
    11'd691 : out <= 24'b11111111111111100000000;
    11'd692 : out <= 24'b11111111111111100000000;
    11'd693 : out <= 24'b11111111111111100000000;
    11'd694 : out <= 24'b00000000000000000000000;
    11'd695 : out <= 24'b00000000000000000000000;
    11'd696 : out <= 24'b00000000000000000000000;
    11'd697 : out <= 24'b00000000000000000000000;
    11'd698 : out <= 24'b0;
    11'd699 : out <= 24'b0;
    11'd700 : out <= 24'b0;
    11'd701 : out <= 24'b0;


// rows 42 to 68
// start rec 26 h = 27 w = 18 ofs = 702
    11'd702 : out <= 24'b00000000000000000000000;
    11'd703 : out <= 24'b00000000000000000000000;
    11'd704 : out <= 24'b00000000000000000000000;
    11'd705 : out <= 24'b00000000000000000000000;
    11'd706 : out <= 24'b00000000000000000000000;
    11'd707 : out <= 24'b00000000000000000000000;
    11'd708 : out <= 24'b01111111111100000000000;
    11'd709 : out <= 24'b01111111111110000000000;
    11'd710 : out <= 24'b01111111111111000000000;
    11'd711 : out <= 24'b00000000001111000000000;
    11'd712 : out <= 24'b00000000000111000000000;
    11'd713 : out <= 24'b00000000000111000000000;
    11'd714 : out <= 24'b00011111111111000000000;
    11'd715 : out <= 24'b01111111111111000000000;
    11'd716 : out <= 24'b11111100011111000000000;
    11'd717 : out <= 24'b11110000001111000000000;
    11'd718 : out <= 24'b11110001111111000000000;
    11'd719 : out <= 24'b11111111111111111000000;
    11'd720 : out <= 24'b01111111111111111000000;
    11'd721 : out <= 24'b00111111100111111000000;
    11'd722 : out <= 24'b00000000000000000000000;
    11'd723 : out <= 24'b00000000000000000000000;
    11'd724 : out <= 24'b00000000000000000000000;
    11'd725 : out <= 24'b00000000000000000000000;
    11'd726 : out <= 24'b00000000000000000000000;
    11'd727 : out <= 24'b00000000000000000000000;
    11'd728 : out <= 24'b0;

// start rec 27 h = 27 w = 20 ofs = 729
    11'd729 : out <= 24'b11111100000000000000000;
    11'd730 : out <= 24'b11111100000000000000000;
    11'd731 : out <= 24'b11111100000000000000000;
    11'd732 : out <= 24'b00011100000000000000000;
    11'd733 : out <= 24'b00011100000000000000000;
    11'd734 : out <= 24'b00011100000000000000000;
    11'd735 : out <= 24'b00011101111111100000000;
    11'd736 : out <= 24'b00011111111111110000000;
    11'd737 : out <= 24'b00011111111111111100000;
    11'd738 : out <= 24'b00011111110011111100000;
    11'd739 : out <= 24'b00011111000000111110000;
    11'd740 : out <= 24'b00011110000000011110000;
    11'd741 : out <= 24'b00011100000000001110000;
    11'd742 : out <= 24'b00011100000000001110000;
    11'd743 : out <= 24'b00011110000000011110000;
    11'd744 : out <= 24'b00011110000000011110000;
    11'd745 : out <= 24'b00011111110011111110000;
    11'd746 : out <= 24'b11111111111111111100000;
    11'd747 : out <= 24'b11111111111111111000000;
    11'd748 : out <= 24'b11111101111111100000000;
    11'd749 : out <= 24'b00000000000000000000000;
    11'd750 : out <= 24'b00000000000000000000000;
    11'd751 : out <= 24'b00000000000000000000000;
    11'd752 : out <= 24'b00000000000000000000000;
    11'd753 : out <= 24'b00000000000000000000000;
    11'd754 : out <= 24'b00000000000000000000000;
    11'd755 : out <= 24'b0;

// start rec 28 h = 27 w = 18 ofs = 756
    11'd756 : out <= 24'b00000000000000000000000;
    11'd757 : out <= 24'b00000000000000000000000;
    11'd758 : out <= 24'b00000000000000000000000;
    11'd759 : out <= 24'b00000000000000000000000;
    11'd760 : out <= 24'b00000000000000000000000;
    11'd761 : out <= 24'b00000000000000000000000;
    11'd762 : out <= 24'b00001111111111110000000;
    11'd763 : out <= 24'b00111111111111110000000;
    11'd764 : out <= 24'b01111111111111110000000;
    11'd765 : out <= 24'b01111110001111110000000;
    11'd766 : out <= 24'b11111000000011110000000;
    11'd767 : out <= 24'b11110000000011110000000;
    11'd768 : out <= 24'b11100000000000000000000;
    11'd769 : out <= 24'b11100000000000000000000;
    11'd770 : out <= 24'b11110000000000000000000;
    11'd771 : out <= 24'b11110000000001111000000;
    11'd772 : out <= 24'b11111110000111111000000;
    11'd773 : out <= 24'b01111111111111111000000;
    11'd774 : out <= 24'b00111111111111110000000;
    11'd775 : out <= 24'b00001111111111100000000;
    11'd776 : out <= 24'b00000000000000000000000;
    11'd777 : out <= 24'b00000000000000000000000;
    11'd778 : out <= 24'b00000000000000000000000;
    11'd779 : out <= 24'b00000000000000000000000;
    11'd780 : out <= 24'b00000000000000000000000;
    11'd781 : out <= 24'b00000000000000000000000;
    11'd782 : out <= 24'b0;

// start rec 29 h = 27 w = 20 ofs = 783
    11'd783 : out <= 24'b00000000001111110000000;
    11'd784 : out <= 24'b00000000001111110000000;
    11'd785 : out <= 24'b00000000001111110000000;
    11'd786 : out <= 24'b00000000000001110000000;
    11'd787 : out <= 24'b00000000000001110000000;
    11'd788 : out <= 24'b00000000000001110000000;
    11'd789 : out <= 24'b00001111111101110000000;
    11'd790 : out <= 24'b00011111111111110000000;
    11'd791 : out <= 24'b01111111111111110000000;
    11'd792 : out <= 24'b01111110011111110000000;
    11'd793 : out <= 24'b11111000000111110000000;
    11'd794 : out <= 24'b11110000000011110000000;
    11'd795 : out <= 24'b11100000000001110000000;
    11'd796 : out <= 24'b11100000000001110000000;
    11'd797 : out <= 24'b11110000000011110000000;
    11'd798 : out <= 24'b11110000000011110000000;
    11'd799 : out <= 24'b11111110011111110000000;
    11'd800 : out <= 24'b01111111111111111110000;
    11'd801 : out <= 24'b00111111111111111110000;
    11'd802 : out <= 24'b00001111111101111110000;
    11'd803 : out <= 24'b00000000000000000000000;
    11'd804 : out <= 24'b00000000000000000000000;
    11'd805 : out <= 24'b00000000000000000000000;
    11'd806 : out <= 24'b00000000000000000000000;
    11'd807 : out <= 24'b00000000000000000000000;
    11'd808 : out <= 24'b00000000000000000000000;
    11'd809 : out <= 24'b0;

// start rec 30 h = 27 w = 18 ofs = 810
    11'd810 : out <= 24'b00000000000000000000000;
    11'd811 : out <= 24'b00000000000000000000000;
    11'd812 : out <= 24'b00000000000000000000000;
    11'd813 : out <= 24'b00000000000000000000000;
    11'd814 : out <= 24'b00000000000000000000000;
    11'd815 : out <= 24'b00000000000000000000000;
    11'd816 : out <= 24'b00001111111110000000000;
    11'd817 : out <= 24'b00011111111111100000000;
    11'd818 : out <= 24'b01111111111111110000000;
    11'd819 : out <= 24'b01111110001111110000000;
    11'd820 : out <= 24'b11111000000011111000000;
    11'd821 : out <= 24'b11110000000001111000000;
    11'd822 : out <= 24'b11111111111111111000000;
    11'd823 : out <= 24'b11111111111111111000000;
    11'd824 : out <= 24'b11110000000000000000000;
    11'd825 : out <= 24'b11111000000000000000000;
    11'd826 : out <= 24'b01111110001111111000000;
    11'd827 : out <= 24'b01111111111111111000000;
    11'd828 : out <= 24'b00111111111111111000000;
    11'd829 : out <= 24'b00001111111111100000000;
    11'd830 : out <= 24'b00000000000000000000000;
    11'd831 : out <= 24'b00000000000000000000000;
    11'd832 : out <= 24'b00000000000000000000000;
    11'd833 : out <= 24'b00000000000000000000000;
    11'd834 : out <= 24'b00000000000000000000000;
    11'd835 : out <= 24'b00000000000000000000000;
    11'd836 : out <= 24'b0;

// start rec 31 h = 27 w = 17 ofs = 837
    11'd837 : out <= 24'b00000011111111110000000;
    11'd838 : out <= 24'b00000111111111110000000;
    11'd839 : out <= 24'b00001111111111110000000;
    11'd840 : out <= 24'b00001111100000000000000;
    11'd841 : out <= 24'b00001110000000000000000;
    11'd842 : out <= 24'b00001110000000000000000;
    11'd843 : out <= 24'b11111111111111000000000;
    11'd844 : out <= 24'b11111111111111000000000;
    11'd845 : out <= 24'b11111111111111000000000;
    11'd846 : out <= 24'b00001110000000000000000;
    11'd847 : out <= 24'b00001110000000000000000;
    11'd848 : out <= 24'b00001110000000000000000;
    11'd849 : out <= 24'b00001110000000000000000;
    11'd850 : out <= 24'b00001110000000000000000;
    11'd851 : out <= 24'b00001110000000000000000;
    11'd852 : out <= 24'b00001110000000000000000;
    11'd853 : out <= 24'b00001110000000000000000;
    11'd854 : out <= 24'b11111111111111000000000;
    11'd855 : out <= 24'b11111111111111000000000;
    11'd856 : out <= 24'b11111111111111000000000;
    11'd857 : out <= 24'b00000000000000000000000;
    11'd858 : out <= 24'b00000000000000000000000;
    11'd859 : out <= 24'b00000000000000000000000;
    11'd860 : out <= 24'b00000000000000000000000;
    11'd861 : out <= 24'b00000000000000000000000;
    11'd862 : out <= 24'b00000000000000000000000;
    11'd863 : out <= 24'b0;

// start rec 32 h = 27 w = 19 ofs = 864
    11'd864 : out <= 24'b00000000000000000000000;
    11'd865 : out <= 24'b00000000000000000000000;
    11'd866 : out <= 24'b00000000000000000000000;
    11'd867 : out <= 24'b00000000000000000000000;
    11'd868 : out <= 24'b00000000000000000000000;
    11'd869 : out <= 24'b00000000000000000000000;
    11'd870 : out <= 24'b00001111111111111100000;
    11'd871 : out <= 24'b00111111111111111100000;
    11'd872 : out <= 24'b01111111111111111100000;
    11'd873 : out <= 24'b01111100011111100000000;
    11'd874 : out <= 24'b11111000001111100000000;
    11'd875 : out <= 24'b11110000000111100000000;
    11'd876 : out <= 24'b11100000000011100000000;
    11'd877 : out <= 24'b11100000000011100000000;
    11'd878 : out <= 24'b11110000000111100000000;
    11'd879 : out <= 24'b11111000001111100000000;
    11'd880 : out <= 24'b01111100011111100000000;
    11'd881 : out <= 24'b01111111111111100000000;
    11'd882 : out <= 24'b00111111111111100000000;
    11'd883 : out <= 24'b00001111111011100000000;
    11'd884 : out <= 24'b00000000000011100000000;
    11'd885 : out <= 24'b00000000000111100000000;
    11'd886 : out <= 24'b00000000001111100000000;
    11'd887 : out <= 24'b00011111111111000000000;
    11'd888 : out <= 24'b00011111111111000000000;
    11'd889 : out <= 24'b00011111111100000000000;
    11'd890 : out <= 24'b0;

// start rec 33 h = 27 w = 19 ofs = 891
    11'd891 : out <= 24'b11111100000000000000000;
    11'd892 : out <= 24'b11111100000000000000000;
    11'd893 : out <= 24'b11111100000000000000000;
    11'd894 : out <= 24'b00011100000000000000000;
    11'd895 : out <= 24'b00011100000000000000000;
    11'd896 : out <= 24'b00011100000000000000000;
    11'd897 : out <= 24'b00011111111111000000000;
    11'd898 : out <= 24'b00011111111111100000000;
    11'd899 : out <= 24'b00011111111111110000000;
    11'd900 : out <= 24'b00011111100111110000000;
    11'd901 : out <= 24'b00011100000011110000000;
    11'd902 : out <= 24'b00011100000001110000000;
    11'd903 : out <= 24'b00011100000001110000000;
    11'd904 : out <= 24'b00011100000001110000000;
    11'd905 : out <= 24'b00011100000001110000000;
    11'd906 : out <= 24'b00011100000001110000000;
    11'd907 : out <= 24'b00011100000001110000000;
    11'd908 : out <= 24'b01111111000111111100000;
    11'd909 : out <= 24'b01111111000111111100000;
    11'd910 : out <= 24'b01111111000111111100000;
    11'd911 : out <= 24'b00000000000000000000000;
    11'd912 : out <= 24'b00000000000000000000000;
    11'd913 : out <= 24'b00000000000000000000000;
    11'd914 : out <= 24'b00000000000000000000000;
    11'd915 : out <= 24'b00000000000000000000000;
    11'd916 : out <= 24'b00000000000000000000000;
    11'd917 : out <= 24'b0;

// start rec 34 h = 27 w = 16 ofs = 918
    11'd918 : out <= 24'b00000011100000000000000;
    11'd919 : out <= 24'b00000011100000000000000;
    11'd920 : out <= 24'b00000011100000000000000;
    11'd921 : out <= 24'b00000000000000000000000;
    11'd922 : out <= 24'b00000000000000000000000;
    11'd923 : out <= 24'b00000000000000000000000;
    11'd924 : out <= 24'b01111111100000000000000;
    11'd925 : out <= 24'b01111111100000000000000;
    11'd926 : out <= 24'b01111111100000000000000;
    11'd927 : out <= 24'b00000011100000000000000;
    11'd928 : out <= 24'b00000011100000000000000;
    11'd929 : out <= 24'b00000011100000000000000;
    11'd930 : out <= 24'b00000011100000000000000;
    11'd931 : out <= 24'b00000011100000000000000;
    11'd932 : out <= 24'b00000011100000000000000;
    11'd933 : out <= 24'b00000011100000000000000;
    11'd934 : out <= 24'b00000011100000000000000;
    11'd935 : out <= 24'b11111111111111100000000;
    11'd936 : out <= 24'b11111111111111100000000;
    11'd937 : out <= 24'b11111111111111100000000;
    11'd938 : out <= 24'b00000000000000000000000;
    11'd939 : out <= 24'b00000000000000000000000;
    11'd940 : out <= 24'b00000000000000000000000;
    11'd941 : out <= 24'b00000000000000000000000;
    11'd942 : out <= 24'b00000000000000000000000;
    11'd943 : out <= 24'b00000000000000000000000;
    11'd944 : out <= 24'b0;

// start rec 35 h = 27 w = 13 ofs = 945
    11'd945 : out <= 24'b00000011100000000000000;
    11'd946 : out <= 24'b00000011100000000000000;
    11'd947 : out <= 24'b00000011100000000000000;
    11'd948 : out <= 24'b00000000000000000000000;
    11'd949 : out <= 24'b00000000000000000000000;
    11'd950 : out <= 24'b00000000000000000000000;
    11'd951 : out <= 24'b11111111111100000000000;
    11'd952 : out <= 24'b11111111111100000000000;
    11'd953 : out <= 24'b11111111111100000000000;
    11'd954 : out <= 24'b00000000011100000000000;
    11'd955 : out <= 24'b00000000011100000000000;
    11'd956 : out <= 24'b00000000011100000000000;
    11'd957 : out <= 24'b00000000011100000000000;
    11'd958 : out <= 24'b00000000011100000000000;
    11'd959 : out <= 24'b00000000011100000000000;
    11'd960 : out <= 24'b00000000011100000000000;
    11'd961 : out <= 24'b00000000011100000000000;
    11'd962 : out <= 24'b00000000011100000000000;
    11'd963 : out <= 24'b00000000011100000000000;
    11'd964 : out <= 24'b00000000011100000000000;
    11'd965 : out <= 24'b00000000011100000000000;
    11'd966 : out <= 24'b00000000111100000000000;
    11'd967 : out <= 24'b00000001111100000000000;
    11'd968 : out <= 24'b11111111111000000000000;
    11'd969 : out <= 24'b11111111111000000000000;
    11'd970 : out <= 24'b11111111100000000000000;
    11'd971 : out <= 24'b0;

// start rec 36 h = 27 w = 18 ofs = 972
    11'd972 : out <= 24'b11111100000000000000000;
    11'd973 : out <= 24'b11111100000000000000000;
    11'd974 : out <= 24'b11111100000000000000000;
    11'd975 : out <= 24'b00011100000000000000000;
    11'd976 : out <= 24'b00011100000000000000000;
    11'd977 : out <= 24'b00011100000000000000000;
    11'd978 : out <= 24'b00011100111111110000000;
    11'd979 : out <= 24'b00011100111111110000000;
    11'd980 : out <= 24'b00011100111111110000000;
    11'd981 : out <= 24'b00011100111111000000000;
    11'd982 : out <= 24'b00011111111110000000000;
    11'd983 : out <= 24'b00011111111000000000000;
    11'd984 : out <= 24'b00011111110000000000000;
    11'd985 : out <= 24'b00011111111000000000000;
    11'd986 : out <= 24'b00011111111100000000000;
    11'd987 : out <= 24'b00011100111110000000000;
    11'd988 : out <= 24'b00011100011111100000000;
    11'd989 : out <= 24'b11111100011111111000000;
    11'd990 : out <= 24'b11111100011111111000000;
    11'd991 : out <= 24'b11111100011111111000000;
    11'd992 : out <= 24'b00000000000000000000000;
    11'd993 : out <= 24'b00000000000000000000000;
    11'd994 : out <= 24'b00000000000000000000000;
    11'd995 : out <= 24'b00000000000000000000000;
    11'd996 : out <= 24'b00000000000000000000000;
    11'd997 : out <= 24'b00000000000000000000000;
    11'd998 : out <= 24'b0;

// start rec 37 h = 27 w = 16 ofs = 999
    11'd999 : out <= 24'b01111111100000000000000;
    11'd1000 : out <= 24'b01111111100000000000000;
    11'd1001 : out <= 24'b01111111100000000000000;
    11'd1002 : out <= 24'b00000011100000000000000;
    11'd1003 : out <= 24'b00000011100000000000000;
    11'd1004 : out <= 24'b00000011100000000000000;
    11'd1005 : out <= 24'b00000011100000000000000;
    11'd1006 : out <= 24'b00000011100000000000000;
    11'd1007 : out <= 24'b00000011100000000000000;
    11'd1008 : out <= 24'b00000011100000000000000;
    11'd1009 : out <= 24'b00000011100000000000000;
    11'd1010 : out <= 24'b00000011100000000000000;
    11'd1011 : out <= 24'b00000011100000000000000;
    11'd1012 : out <= 24'b00000011100000000000000;
    11'd1013 : out <= 24'b00000011100000000000000;
    11'd1014 : out <= 24'b00000011100000000000000;
    11'd1015 : out <= 24'b00000011100000000000000;
    11'd1016 : out <= 24'b11111111111111100000000;
    11'd1017 : out <= 24'b11111111111111100000000;
    11'd1018 : out <= 24'b11111111111111100000000;
    11'd1019 : out <= 24'b00000000000000000000000;
    11'd1020 : out <= 24'b00000000000000000000000;
    11'd1021 : out <= 24'b00000000000000000000000;
    11'd1022 : out <= 24'b00000000000000000000000;
    11'd1023 : out <= 24'b00000000000000000000000;
    11'd1024 : out <= 24'b00000000000000000000000;
    11'd1025 : out <= 24'b0;

// start rec 38 h = 27 w = 22 ofs = 1026
    11'd1026 : out <= 24'b00000000000000000000000;
    11'd1027 : out <= 24'b00000000000000000000000;
    11'd1028 : out <= 24'b00000000000000000000000;
    11'd1029 : out <= 24'b00000000000000000000000;
    11'd1030 : out <= 24'b00000000000000000000000;
    11'd1031 : out <= 24'b00000000000000000000000;
    11'd1032 : out <= 24'b11111011110011111100000;
    11'd1033 : out <= 24'b11111111111111111110000;
    11'd1034 : out <= 24'b11111111111111111110000;
    11'd1035 : out <= 24'b00111110111111011110000;
    11'd1036 : out <= 24'b00111100011110001110000;
    11'd1037 : out <= 24'b00111000011100001110000;
    11'd1038 : out <= 24'b00111000011100001110000;
    11'd1039 : out <= 24'b00111000011100001110000;
    11'd1040 : out <= 24'b00111000011100001110000;
    11'd1041 : out <= 24'b00111000011100001110000;
    11'd1042 : out <= 24'b00111000011100001110000;
    11'd1043 : out <= 24'b11111110011111001111100;
    11'd1044 : out <= 24'b11111110011111001111100;
    11'd1045 : out <= 24'b11111110011111001111100;
    11'd1046 : out <= 24'b00000000000000000000000;
    11'd1047 : out <= 24'b00000000000000000000000;
    11'd1048 : out <= 24'b00000000000000000000000;
    11'd1049 : out <= 24'b00000000000000000000000;
    11'd1050 : out <= 24'b00000000000000000000000;
    11'd1051 : out <= 24'b00000000000000000000000;
    11'd1052 : out <= 24'b0;

// start rec 39 h = 27 w = 18 ofs = 1053
    11'd1053 : out <= 24'b00000000000000000000000;
    11'd1054 : out <= 24'b00000000000000000000000;
    11'd1055 : out <= 24'b00000000000000000000000;
    11'd1056 : out <= 24'b00000000000000000000000;
    11'd1057 : out <= 24'b00000000000000000000000;
    11'd1058 : out <= 24'b00000000000000000000000;
    11'd1059 : out <= 24'b11111111111110000000000;
    11'd1060 : out <= 24'b11111111111111000000000;
    11'd1061 : out <= 24'b11111111111111100000000;
    11'd1062 : out <= 24'b00111111001111100000000;
    11'd1063 : out <= 24'b00111000000011100000000;
    11'd1064 : out <= 24'b00111000000011100000000;
    11'd1065 : out <= 24'b00111000000011100000000;
    11'd1066 : out <= 24'b00111000000011100000000;
    11'd1067 : out <= 24'b00111000000011100000000;
    11'd1068 : out <= 24'b00111000000011100000000;
    11'd1069 : out <= 24'b00111000000011100000000;
    11'd1070 : out <= 24'b11111110001111111000000;
    11'd1071 : out <= 24'b11111110001111111000000;
    11'd1072 : out <= 24'b11111110001111111000000;
    11'd1073 : out <= 24'b00000000000000000000000;
    11'd1074 : out <= 24'b00000000000000000000000;
    11'd1075 : out <= 24'b00000000000000000000000;
    11'd1076 : out <= 24'b00000000000000000000000;
    11'd1077 : out <= 24'b00000000000000000000000;
    11'd1078 : out <= 24'b00000000000000000000000;
    11'd1079 : out <= 24'b0;

// start rec 40 h = 27 w = 18 ofs = 1080
    11'd1080 : out <= 24'b00000000000000000000000;
    11'd1081 : out <= 24'b00000000000000000000000;
    11'd1082 : out <= 24'b00000000000000000000000;
    11'd1083 : out <= 24'b00000000000000000000000;
    11'd1084 : out <= 24'b00000000000000000000000;
    11'd1085 : out <= 24'b00000000000000000000000;
    11'd1086 : out <= 24'b00001111111110000000000;
    11'd1087 : out <= 24'b00011111111111000000000;
    11'd1088 : out <= 24'b00111111111111100000000;
    11'd1089 : out <= 24'b01111110001111110000000;
    11'd1090 : out <= 24'b11111000000011111000000;
    11'd1091 : out <= 24'b11110000000001111000000;
    11'd1092 : out <= 24'b11100000000000111000000;
    11'd1093 : out <= 24'b11100000000000111000000;
    11'd1094 : out <= 24'b11110000000001111000000;
    11'd1095 : out <= 24'b11111000000011111000000;
    11'd1096 : out <= 24'b01111110001111110000000;
    11'd1097 : out <= 24'b01111111111111110000000;
    11'd1098 : out <= 24'b00111111111111100000000;
    11'd1099 : out <= 24'b00001111111110000000000;
    11'd1100 : out <= 24'b00000000000000000000000;
    11'd1101 : out <= 24'b00000000000000000000000;
    11'd1102 : out <= 24'b00000000000000000000000;
    11'd1103 : out <= 24'b00000000000000000000000;
    11'd1104 : out <= 24'b00000000000000000000000;
    11'd1105 : out <= 24'b00000000000000000000000;
    11'd1106 : out <= 24'b0;

// start rec 41 h = 27 w = 20 ofs = 1107
    11'd1107 : out <= 24'b00000000000000000000000;
    11'd1108 : out <= 24'b00000000000000000000000;
    11'd1109 : out <= 24'b00000000000000000000000;
    11'd1110 : out <= 24'b00000000000000000000000;
    11'd1111 : out <= 24'b00000000000000000000000;
    11'd1112 : out <= 24'b00000000000000000000000;
    11'd1113 : out <= 24'b11111111111111100000000;
    11'd1114 : out <= 24'b11111111111111110000000;
    11'd1115 : out <= 24'b11111111111111111000000;
    11'd1116 : out <= 24'b00011111110011111100000;
    11'd1117 : out <= 24'b00011111000000111110000;
    11'd1118 : out <= 24'b00011110000000011110000;
    11'd1119 : out <= 24'b00011110000000011110000;
    11'd1120 : out <= 24'b00011100000000001110000;
    11'd1121 : out <= 24'b00011110000000011110000;
    11'd1122 : out <= 24'b00011111000000111110000;
    11'd1123 : out <= 24'b00011111110011111100000;
    11'd1124 : out <= 24'b00011111111111111100000;
    11'd1125 : out <= 24'b00011111111111111000000;
    11'd1126 : out <= 24'b00011101111111100000000;
    11'd1127 : out <= 24'b00011100000000000000000;
    11'd1128 : out <= 24'b00011100000000000000000;
    11'd1129 : out <= 24'b00011100000000000000000;
    11'd1130 : out <= 24'b11111111110000000000000;
    11'd1131 : out <= 24'b11111111110000000000000;
    11'd1132 : out <= 24'b11111111110000000000000;
    11'd1133 : out <= 24'b0;

// start rec 42 h = 27 w = 20 ofs = 1134
    11'd1134 : out <= 24'b00000000000000000000000;
    11'd1135 : out <= 24'b00000000000000000000000;
    11'd1136 : out <= 24'b00000000000000000000000;
    11'd1137 : out <= 24'b00000000000000000000000;
    11'd1138 : out <= 24'b00000000000000000000000;
    11'd1139 : out <= 24'b00000000000000000000000;
    11'd1140 : out <= 24'b00001111111111111110000;
    11'd1141 : out <= 24'b00011111111111111110000;
    11'd1142 : out <= 24'b00111111111111111110000;
    11'd1143 : out <= 24'b01111110011111110000000;
    11'd1144 : out <= 24'b11111000000111110000000;
    11'd1145 : out <= 24'b11110000000011110000000;
    11'd1146 : out <= 24'b11110000000011110000000;
    11'd1147 : out <= 24'b11100000000001110000000;
    11'd1148 : out <= 24'b11110000000011110000000;
    11'd1149 : out <= 24'b11111000000111110000000;
    11'd1150 : out <= 24'b01111110011111110000000;
    11'd1151 : out <= 24'b01111111111111110000000;
    11'd1152 : out <= 24'b00111111111111110000000;
    11'd1153 : out <= 24'b00001111111101110000000;
    11'd1154 : out <= 24'b00000000000001110000000;
    11'd1155 : out <= 24'b00000000000001110000000;
    11'd1156 : out <= 24'b00000000000001110000000;
    11'd1157 : out <= 24'b00000000011111111110000;
    11'd1158 : out <= 24'b00000000011111111110000;
    11'd1159 : out <= 24'b00000000011111111110000;
    11'd1160 : out <= 24'b0;

// start rec 43 h = 27 w = 17 ofs = 1161
    11'd1161 : out <= 24'b00000000000000000000000;
    11'd1162 : out <= 24'b00000000000000000000000;
    11'd1163 : out <= 24'b00000000000000000000000;
    11'd1164 : out <= 24'b00000000000000000000000;
    11'd1165 : out <= 24'b00000000000000000000000;
    11'd1166 : out <= 24'b00000000000000000000000;
    11'd1167 : out <= 24'b01111110001111100000000;
    11'd1168 : out <= 24'b01111110111111110000000;
    11'd1169 : out <= 24'b01111111111111110000000;
    11'd1170 : out <= 24'b00001111111101110000000;
    11'd1171 : out <= 24'b00001111110000000000000;
    11'd1172 : out <= 24'b00001111100000000000000;
    11'd1173 : out <= 24'b00001110000000000000000;
    11'd1174 : out <= 24'b00001110000000000000000;
    11'd1175 : out <= 24'b00001110000000000000000;
    11'd1176 : out <= 24'b00001110000000000000000;
    11'd1177 : out <= 24'b00001110000000000000000;
    11'd1178 : out <= 24'b11111111111111000000000;
    11'd1179 : out <= 24'b11111111111111000000000;
    11'd1180 : out <= 24'b11111111111111000000000;
    11'd1181 : out <= 24'b00000000000000000000000;
    11'd1182 : out <= 24'b00000000000000000000000;
    11'd1183 : out <= 24'b00000000000000000000000;
    11'd1184 : out <= 24'b00000000000000000000000;
    11'd1185 : out <= 24'b00000000000000000000000;
    11'd1186 : out <= 24'b00000000000000000000000;
    11'd1187 : out <= 24'b0;

// start rec 44 h = 27 w = 16 ofs = 1188
    11'd1188 : out <= 24'b00000000000000000000000;
    11'd1189 : out <= 24'b00000000000000000000000;
    11'd1190 : out <= 24'b00000000000000000000000;
    11'd1191 : out <= 24'b00000000000000000000000;
    11'd1192 : out <= 24'b00000000000000000000000;
    11'd1193 : out <= 24'b00000000000000000000000;
    11'd1194 : out <= 24'b00011111111111000000000;
    11'd1195 : out <= 24'b00111111111111000000000;
    11'd1196 : out <= 24'b01111111111111000000000;
    11'd1197 : out <= 24'b01111100011111000000000;
    11'd1198 : out <= 24'b01111000000111000000000;
    11'd1199 : out <= 24'b01111111111000000000000;
    11'd1200 : out <= 24'b00111111111111000000000;
    11'd1201 : out <= 24'b00011111111111100000000;
    11'd1202 : out <= 24'b00000001111111100000000;
    11'd1203 : out <= 24'b11110000000011100000000;
    11'd1204 : out <= 24'b11111100001111100000000;
    11'd1205 : out <= 24'b11111111111111100000000;
    11'd1206 : out <= 24'b11111111111111000000000;
    11'd1207 : out <= 24'b11111111111100000000000;
    11'd1208 : out <= 24'b00000000000000000000000;
    11'd1209 : out <= 24'b00000000000000000000000;
    11'd1210 : out <= 24'b00000000000000000000000;
    11'd1211 : out <= 24'b00000000000000000000000;
    11'd1212 : out <= 24'b00000000000000000000000;
    11'd1213 : out <= 24'b00000000000000000000000;
    11'd1214 : out <= 24'b0;

// start rec 45 h = 27 w = 17 ofs = 1215
    11'd1215 : out <= 24'b00000000000000000000000;
    11'd1216 : out <= 24'b00011100000000000000000;
    11'd1217 : out <= 24'b00011100000000000000000;
    11'd1218 : out <= 24'b00011100000000000000000;
    11'd1219 : out <= 24'b00011100000000000000000;
    11'd1220 : out <= 24'b00011100000000000000000;
    11'd1221 : out <= 24'b11111111111111000000000;
    11'd1222 : out <= 24'b11111111111111000000000;
    11'd1223 : out <= 24'b11111111111111000000000;
    11'd1224 : out <= 24'b00011100000000000000000;
    11'd1225 : out <= 24'b00011100000000000000000;
    11'd1226 : out <= 24'b00011100000000000000000;
    11'd1227 : out <= 24'b00011100000000000000000;
    11'd1228 : out <= 24'b00011100000000000000000;
    11'd1229 : out <= 24'b00011100000000000000000;
    11'd1230 : out <= 24'b00011100000000000000000;
    11'd1231 : out <= 24'b00011110000111110000000;
    11'd1232 : out <= 24'b00011111111111110000000;
    11'd1233 : out <= 24'b00001111111111110000000;
    11'd1234 : out <= 24'b00000111111111000000000;
    11'd1235 : out <= 24'b00000000000000000000000;
    11'd1236 : out <= 24'b00000000000000000000000;
    11'd1237 : out <= 24'b00000000000000000000000;
    11'd1238 : out <= 24'b00000000000000000000000;
    11'd1239 : out <= 24'b00000000000000000000000;
    11'd1240 : out <= 24'b00000000000000000000000;
    11'd1241 : out <= 24'b0;

// start rec 46 h = 27 w = 19 ofs = 1242
    11'd1242 : out <= 24'b00000000000000000000000;
    11'd1243 : out <= 24'b00000000000000000000000;
    11'd1244 : out <= 24'b00000000000000000000000;
    11'd1245 : out <= 24'b00000000000000000000000;
    11'd1246 : out <= 24'b00000000000000000000000;
    11'd1247 : out <= 24'b00000000000000000000000;
    11'd1248 : out <= 24'b11111100001111110000000;
    11'd1249 : out <= 24'b11111100001111110000000;
    11'd1250 : out <= 24'b11111100001111110000000;
    11'd1251 : out <= 24'b00011100000001110000000;
    11'd1252 : out <= 24'b00011100000001110000000;
    11'd1253 : out <= 24'b00011100000001110000000;
    11'd1254 : out <= 24'b00011100000001110000000;
    11'd1255 : out <= 24'b00011100000001110000000;
    11'd1256 : out <= 24'b00011100000001110000000;
    11'd1257 : out <= 24'b00011100000011110000000;
    11'd1258 : out <= 24'b00011110011111110000000;
    11'd1259 : out <= 24'b00011111111111111100000;
    11'd1260 : out <= 24'b00001111111111111100000;
    11'd1261 : out <= 24'b00000111111111111100000;
    11'd1262 : out <= 24'b00000000000000000000000;
    11'd1263 : out <= 24'b00000000000000000000000;
    11'd1264 : out <= 24'b00000000000000000000000;
    11'd1265 : out <= 24'b00000000000000000000000;
    11'd1266 : out <= 24'b00000000000000000000000;
    11'd1267 : out <= 24'b00000000000000000000000;
    11'd1268 : out <= 24'b0;

// start rec 47 h = 27 w = 19 ofs = 1269
    11'd1269 : out <= 24'b00000000000000000000000;
    11'd1270 : out <= 24'b00000000000000000000000;
    11'd1271 : out <= 24'b00000000000000000000000;
    11'd1272 : out <= 24'b00000000000000000000000;
    11'd1273 : out <= 24'b00000000000000000000000;
    11'd1274 : out <= 24'b00000000000000000000000;
    11'd1275 : out <= 24'b11111110001111111100000;
    11'd1276 : out <= 24'b11111110001111111100000;
    11'd1277 : out <= 24'b11111110001111111100000;
    11'd1278 : out <= 24'b00111100000111100000000;
    11'd1279 : out <= 24'b00111100000111100000000;
    11'd1280 : out <= 24'b00011100000111000000000;
    11'd1281 : out <= 24'b00011110001111000000000;
    11'd1282 : out <= 24'b00011110001111000000000;
    11'd1283 : out <= 24'b00001111011110000000000;
    11'd1284 : out <= 24'b00001111011110000000000;
    11'd1285 : out <= 24'b00000111111100000000000;
    11'd1286 : out <= 24'b00000111111100000000000;
    11'd1287 : out <= 24'b00000111111100000000000;
    11'd1288 : out <= 24'b00000011111000000000000;
    11'd1289 : out <= 24'b00000000000000000000000;
    11'd1290 : out <= 24'b00000000000000000000000;
    11'd1291 : out <= 24'b00000000000000000000000;
    11'd1292 : out <= 24'b00000000000000000000000;
    11'd1293 : out <= 24'b00000000000000000000000;
    11'd1294 : out <= 24'b00000000000000000000000;
    11'd1295 : out <= 24'b0;

// start rec 48 h = 27 w = 20 ofs = 1296
    11'd1296 : out <= 24'b00000000000000000000000;
    11'd1297 : out <= 24'b00000000000000000000000;
    11'd1298 : out <= 24'b00000000000000000000000;
    11'd1299 : out <= 24'b00000000000000000000000;
    11'd1300 : out <= 24'b00000000000000000000000;
    11'd1301 : out <= 24'b00000000000000000000000;
    11'd1302 : out <= 24'b11111110000011111110000;
    11'd1303 : out <= 24'b11111110000011111110000;
    11'd1304 : out <= 24'b11111110000011111110000;
    11'd1305 : out <= 24'b00111000111000111000000;
    11'd1306 : out <= 24'b00111001111100111000000;
    11'd1307 : out <= 24'b00111101111101111000000;
    11'd1308 : out <= 24'b00011101111101110000000;
    11'd1309 : out <= 24'b00011111111111110000000;
    11'd1310 : out <= 24'b00011111101111110000000;
    11'd1311 : out <= 24'b00011111101111110000000;
    11'd1312 : out <= 24'b00001111001111100000000;
    11'd1313 : out <= 24'b00001111000111100000000;
    11'd1314 : out <= 24'b00001111000111100000000;
    11'd1315 : out <= 24'b00001110000111100000000;
    11'd1316 : out <= 24'b00000000000000000000000;
    11'd1317 : out <= 24'b00000000000000000000000;
    11'd1318 : out <= 24'b00000000000000000000000;
    11'd1319 : out <= 24'b00000000000000000000000;
    11'd1320 : out <= 24'b00000000000000000000000;
    11'd1321 : out <= 24'b00000000000000000000000;
    11'd1322 : out <= 24'b0;

// start rec 49 h = 27 w = 18 ofs = 1323
    11'd1323 : out <= 24'b00000000000000000000000;
    11'd1324 : out <= 24'b00000000000000000000000;
    11'd1325 : out <= 24'b00000000000000000000000;
    11'd1326 : out <= 24'b00000000000000000000000;
    11'd1327 : out <= 24'b00000000000000000000000;
    11'd1328 : out <= 24'b00000000000000000000000;
    11'd1329 : out <= 24'b01111111011111110000000;
    11'd1330 : out <= 24'b01111111011111110000000;
    11'd1331 : out <= 24'b01111111011111110000000;
    11'd1332 : out <= 24'b00001111011110000000000;
    11'd1333 : out <= 24'b00000111111100000000000;
    11'd1334 : out <= 24'b00000111111000000000000;
    11'd1335 : out <= 24'b00000011111000000000000;
    11'd1336 : out <= 24'b00000011111000000000000;
    11'd1337 : out <= 24'b00000111111100000000000;
    11'd1338 : out <= 24'b00001111011110000000000;
    11'd1339 : out <= 24'b00011110001111000000000;
    11'd1340 : out <= 24'b11111110001111111000000;
    11'd1341 : out <= 24'b11111110001111111000000;
    11'd1342 : out <= 24'b11111110001111111000000;
    11'd1343 : out <= 24'b00000000000000000000000;
    11'd1344 : out <= 24'b00000000000000000000000;
    11'd1345 : out <= 24'b00000000000000000000000;
    11'd1346 : out <= 24'b00000000000000000000000;
    11'd1347 : out <= 24'b00000000000000000000000;
    11'd1348 : out <= 24'b00000000000000000000000;
    11'd1349 : out <= 24'b0;

// start rec 50 h = 27 w = 19 ofs = 1350
    11'd1350 : out <= 24'b00000000000000000000000;
    11'd1351 : out <= 24'b00000000000000000000000;
    11'd1352 : out <= 24'b00000000000000000000000;
    11'd1353 : out <= 24'b00000000000000000000000;
    11'd1354 : out <= 24'b00000000000000000000000;
    11'd1355 : out <= 24'b00000000000000000000000;
    11'd1356 : out <= 24'b11111110000111111100000;
    11'd1357 : out <= 24'b11111110000111111100000;
    11'd1358 : out <= 24'b11111110000111111100000;
    11'd1359 : out <= 24'b00111100000011110000000;
    11'd1360 : out <= 24'b00111100000011110000000;
    11'd1361 : out <= 24'b00011110000111100000000;
    11'd1362 : out <= 24'b00001110000111100000000;
    11'd1363 : out <= 24'b00001111001111000000000;
    11'd1364 : out <= 24'b00000111101111000000000;
    11'd1365 : out <= 24'b00000111111110000000000;
    11'd1366 : out <= 24'b00000011111110000000000;
    11'd1367 : out <= 24'b00000011111100000000000;
    11'd1368 : out <= 24'b00000001111100000000000;
    11'd1369 : out <= 24'b00000001111000000000000;
    11'd1370 : out <= 24'b00000011111000000000000;
    11'd1371 : out <= 24'b00000011110000000000000;
    11'd1372 : out <= 24'b00000011110000000000000;
    11'd1373 : out <= 24'b01111111111100000000000;
    11'd1374 : out <= 24'b01111111111100000000000;
    11'd1375 : out <= 24'b01111111111100000000000;
    11'd1376 : out <= 24'b0;

// start rec 51 h = 27 w = 14 ofs = 1377
    11'd1377 : out <= 24'b00000000000000000000000;
    11'd1378 : out <= 24'b00000000000000000000000;
    11'd1379 : out <= 24'b00000000000000000000000;
    11'd1380 : out <= 24'b00000000000000000000000;
    11'd1381 : out <= 24'b00000000000000000000000;
    11'd1382 : out <= 24'b00000000000000000000000;
    11'd1383 : out <= 24'b11111111111110000000000;
    11'd1384 : out <= 24'b11111111111110000000000;
    11'd1385 : out <= 24'b11111111111110000000000;
    11'd1386 : out <= 24'b11100000111110000000000;
    11'd1387 : out <= 24'b11100001111000000000000;
    11'd1388 : out <= 24'b00000011110000000000000;
    11'd1389 : out <= 24'b00000111100000000000000;
    11'd1390 : out <= 24'b00001111000000000000000;
    11'd1391 : out <= 24'b00011110000000000000000;
    11'd1392 : out <= 24'b00111100001110000000000;
    11'd1393 : out <= 24'b11111000001110000000000;
    11'd1394 : out <= 24'b11111111111110000000000;
    11'd1395 : out <= 24'b11111111111110000000000;
    11'd1396 : out <= 24'b11111111111110000000000;
    11'd1397 : out <= 24'b00000000000000000000000;
    11'd1398 : out <= 24'b00000000000000000000000;
    11'd1399 : out <= 24'b00000000000000000000000;
    11'd1400 : out <= 24'b00000000000000000000000;
    11'd1401 : out <= 24'b00000000000000000000000;
    11'd1402 : out <= 24'b00000000000000000000000;
    11'd1403 : out <= 24'b0;


// rows 76 to 102
// start rec 52 h = 27 w = 15 ofs = 1404
    11'd1404 : out <= 24'b00000000000000000000000;
    11'd1405 : out <= 24'b00000000000000000000000;
    11'd1406 : out <= 24'b00001111110000000000000;
    11'd1407 : out <= 24'b00111111111100000000000;
    11'd1408 : out <= 24'b01111111111100000000000;
    11'd1409 : out <= 24'b01111100111110000000000;
    11'd1410 : out <= 24'b11111000011111000000000;
    11'd1411 : out <= 24'b11110000001111000000000;
    11'd1412 : out <= 24'b11110000001111000000000;
    11'd1413 : out <= 24'b11100000000111000000000;
    11'd1414 : out <= 24'b11100000000111000000000;
    11'd1415 : out <= 24'b11100000000111000000000;
    11'd1416 : out <= 24'b11100000000111000000000;
    11'd1417 : out <= 24'b11100000000111000000000;
    11'd1418 : out <= 24'b11100000000111000000000;
    11'd1419 : out <= 24'b11110000001111000000000;
    11'd1420 : out <= 24'b11110000001111000000000;
    11'd1421 : out <= 24'b11111000011111000000000;
    11'd1422 : out <= 24'b01111100111110000000000;
    11'd1423 : out <= 24'b00111111111110000000000;
    11'd1424 : out <= 24'b00111111111100000000000;
    11'd1425 : out <= 24'b00011111110000000000000;
    11'd1426 : out <= 24'b00000000000000000000000;
    11'd1427 : out <= 24'b00000000000000000000000;
    11'd1428 : out <= 24'b00000000000000000000000;
    11'd1429 : out <= 24'b00000000000000000000000;
    11'd1430 : out <= 24'b0;

// start rec 53 h = 27 w = 14 ofs = 1431
    11'd1431 : out <= 24'b00000000000000000000000;
    11'd1432 : out <= 24'b00000000000000000000000;
    11'd1433 : out <= 24'b00000111000000000000000;
    11'd1434 : out <= 24'b01111111000000000000000;
    11'd1435 : out <= 24'b11111111000000000000000;
    11'd1436 : out <= 24'b11111111000000000000000;
    11'd1437 : out <= 24'b11111111000000000000000;
    11'd1438 : out <= 24'b00000111000000000000000;
    11'd1439 : out <= 24'b00000111000000000000000;
    11'd1440 : out <= 24'b00000111000000000000000;
    11'd1441 : out <= 24'b00000111000000000000000;
    11'd1442 : out <= 24'b00000111000000000000000;
    11'd1443 : out <= 24'b00000111000000000000000;
    11'd1444 : out <= 24'b00000111000000000000000;
    11'd1445 : out <= 24'b00000111000000000000000;
    11'd1446 : out <= 24'b00000111000000000000000;
    11'd1447 : out <= 24'b00000111000000000000000;
    11'd1448 : out <= 24'b00000111000000000000000;
    11'd1449 : out <= 24'b00000111000000000000000;
    11'd1450 : out <= 24'b11111111111110000000000;
    11'd1451 : out <= 24'b11111111111110000000000;
    11'd1452 : out <= 24'b11111111111110000000000;
    11'd1453 : out <= 24'b00000000000000000000000;
    11'd1454 : out <= 24'b00000000000000000000000;
    11'd1455 : out <= 24'b00000000000000000000000;
    11'd1456 : out <= 24'b00000000000000000000000;
    11'd1457 : out <= 24'b0;

// start rec 54 h = 27 w = 15 ofs = 1458
    11'd1458 : out <= 24'b00000000000000000000000;
    11'd1459 : out <= 24'b00000000000000000000000;
    11'd1460 : out <= 24'b00001111111000000000000;
    11'd1461 : out <= 24'b00011111111100000000000;
    11'd1462 : out <= 24'b00111111111110000000000;
    11'd1463 : out <= 24'b01111110111111000000000;
    11'd1464 : out <= 24'b01111000001111000000000;
    11'd1465 : out <= 24'b01110000000111000000000;
    11'd1466 : out <= 24'b01110000000111000000000;
    11'd1467 : out <= 24'b00000000001111000000000;
    11'd1468 : out <= 24'b00000000011111000000000;
    11'd1469 : out <= 24'b00000000111110000000000;
    11'd1470 : out <= 24'b00000001111100000000000;
    11'd1471 : out <= 24'b00000011111000000000000;
    11'd1472 : out <= 24'b00000111110000000000000;
    11'd1473 : out <= 24'b00001111000000000000000;
    11'd1474 : out <= 24'b00111110000000000000000;
    11'd1475 : out <= 24'b01111100000000000000000;
    11'd1476 : out <= 24'b11110000000000000000000;
    11'd1477 : out <= 24'b11111111111111000000000;
    11'd1478 : out <= 24'b11111111111111000000000;
    11'd1479 : out <= 24'b11111111111111000000000;
    11'd1480 : out <= 24'b00000000000000000000000;
    11'd1481 : out <= 24'b00000000000000000000000;
    11'd1482 : out <= 24'b00000000000000000000000;
    11'd1483 : out <= 24'b00000000000000000000000;
    11'd1484 : out <= 24'b0;

// start rec 55 h = 27 w = 16 ofs = 1485
    11'd1485 : out <= 24'b00000000000000000000000;
    11'd1486 : out <= 24'b00000000000000000000000;
    11'd1487 : out <= 24'b00011111111000000000000;
    11'd1488 : out <= 24'b00111111111110000000000;
    11'd1489 : out <= 24'b01111111111110000000000;
    11'd1490 : out <= 24'b01111100011111000000000;
    11'd1491 : out <= 24'b01110000001111000000000;
    11'd1492 : out <= 24'b00000000000111000000000;
    11'd1493 : out <= 24'b00000000001111000000000;
    11'd1494 : out <= 24'b00000000011111000000000;
    11'd1495 : out <= 24'b00000111111110000000000;
    11'd1496 : out <= 24'b00000111111110000000000;
    11'd1497 : out <= 24'b00000111111111000000000;
    11'd1498 : out <= 24'b00000000111111100000000;
    11'd1499 : out <= 24'b00000000000111100000000;
    11'd1500 : out <= 24'b00000000000111100000000;
    11'd1501 : out <= 24'b00000000000011100000000;
    11'd1502 : out <= 24'b00000000000111100000000;
    11'd1503 : out <= 24'b11110000011111100000000;
    11'd1504 : out <= 24'b11111111111111000000000;
    11'd1505 : out <= 24'b11111111111110000000000;
    11'd1506 : out <= 24'b01111111111100000000000;
    11'd1507 : out <= 24'b00000000000000000000000;
    11'd1508 : out <= 24'b00000000000000000000000;
    11'd1509 : out <= 24'b00000000000000000000000;
    11'd1510 : out <= 24'b00000000000000000000000;
    11'd1511 : out <= 24'b0;

// start rec 56 h = 27 w = 15 ofs = 1512
    11'd1512 : out <= 24'b00000000000000000000000;
    11'd1513 : out <= 24'b00000000000000000000000;
    11'd1514 : out <= 24'b00000001111100000000000;
    11'd1515 : out <= 24'b00000001111100000000000;
    11'd1516 : out <= 24'b00000011111100000000000;
    11'd1517 : out <= 24'b00000111111100000000000;
    11'd1518 : out <= 24'b00000111111100000000000;
    11'd1519 : out <= 24'b00001111011100000000000;
    11'd1520 : out <= 24'b00011110011100000000000;
    11'd1521 : out <= 24'b00011110011100000000000;
    11'd1522 : out <= 24'b00111100011100000000000;
    11'd1523 : out <= 24'b01111100011100000000000;
    11'd1524 : out <= 24'b01111000011100000000000;
    11'd1525 : out <= 24'b11110000011100000000000;
    11'd1526 : out <= 24'b11111111111111000000000;
    11'd1527 : out <= 24'b11111111111111000000000;
    11'd1528 : out <= 24'b11111111111111000000000;
    11'd1529 : out <= 24'b00000000011100000000000;
    11'd1530 : out <= 24'b00000000011100000000000;
    11'd1531 : out <= 24'b00000011111111000000000;
    11'd1532 : out <= 24'b00000011111111000000000;
    11'd1533 : out <= 24'b00000011111111000000000;
    11'd1534 : out <= 24'b00000000000000000000000;
    11'd1535 : out <= 24'b00000000000000000000000;
    11'd1536 : out <= 24'b00000000000000000000000;
    11'd1537 : out <= 24'b00000000000000000000000;
    11'd1538 : out <= 24'b0;

// start rec 57 h = 27 w = 16 ofs = 1539
    11'd1539 : out <= 24'b00000000000000000000000;
    11'd1540 : out <= 24'b00000000000000000000000;
    11'd1541 : out <= 24'b00111111111111000000000;
    11'd1542 : out <= 24'b00111111111111000000000;
    11'd1543 : out <= 24'b00111111111111000000000;
    11'd1544 : out <= 24'b00111000000000000000000;
    11'd1545 : out <= 24'b00111000000000000000000;
    11'd1546 : out <= 24'b00111000000000000000000;
    11'd1547 : out <= 24'b00111111111100000000000;
    11'd1548 : out <= 24'b00111111111110000000000;
    11'd1549 : out <= 24'b00111111111111000000000;
    11'd1550 : out <= 24'b00111111011111100000000;
    11'd1551 : out <= 24'b00111000000111100000000;
    11'd1552 : out <= 24'b00000000000111100000000;
    11'd1553 : out <= 24'b00000000000011100000000;
    11'd1554 : out <= 24'b00000000000011100000000;
    11'd1555 : out <= 24'b00000000000111100000000;
    11'd1556 : out <= 24'b11100000000111100000000;
    11'd1557 : out <= 24'b11111000011111100000000;
    11'd1558 : out <= 24'b11111111111111000000000;
    11'd1559 : out <= 24'b01111111111110000000000;
    11'd1560 : out <= 24'b00111111111100000000000;
    11'd1561 : out <= 24'b00000000000000000000000;
    11'd1562 : out <= 24'b00000000000000000000000;
    11'd1563 : out <= 24'b00000000000000000000000;
    11'd1564 : out <= 24'b00000000000000000000000;
    11'd1565 : out <= 24'b0;

// start rec 58 h = 27 w = 15 ofs = 1566
    11'd1566 : out <= 24'b00000000000000000000000;
    11'd1567 : out <= 24'b00000000000000000000000;
    11'd1568 : out <= 24'b00000011111110000000000;
    11'd1569 : out <= 24'b00001111111111000000000;
    11'd1570 : out <= 24'b00011111111111000000000;
    11'd1571 : out <= 24'b00111111100111000000000;
    11'd1572 : out <= 24'b01111110000000000000000;
    11'd1573 : out <= 24'b01111000000000000000000;
    11'd1574 : out <= 24'b11110000000000000000000;
    11'd1575 : out <= 24'b11111111111000000000000;
    11'd1576 : out <= 24'b11111111111100000000000;
    11'd1577 : out <= 24'b11111111111110000000000;
    11'd1578 : out <= 24'b11111110111111000000000;
    11'd1579 : out <= 24'b11111000001111000000000;
    11'd1580 : out <= 24'b11110000001111000000000;
    11'd1581 : out <= 24'b11110000000111000000000;
    11'd1582 : out <= 24'b11110000000111000000000;
    11'd1583 : out <= 24'b11110000001111000000000;
    11'd1584 : out <= 24'b01111100111111000000000;
    11'd1585 : out <= 24'b01111111111110000000000;
    11'd1586 : out <= 24'b00111111111110000000000;
    11'd1587 : out <= 24'b00001111111000000000000;
    11'd1588 : out <= 24'b00000000000000000000000;
    11'd1589 : out <= 24'b00000000000000000000000;
    11'd1590 : out <= 24'b00000000000000000000000;
    11'd1591 : out <= 24'b00000000000000000000000;
    11'd1592 : out <= 24'b0;

// start rec 59 h = 27 w = 14 ofs = 1593
    11'd1593 : out <= 24'b00000000000000000000000;
    11'd1594 : out <= 24'b00000000000000000000000;
    11'd1595 : out <= 24'b11111111111110000000000;
    11'd1596 : out <= 24'b11111111111110000000000;
    11'd1597 : out <= 24'b11111111111110000000000;
    11'd1598 : out <= 24'b11100000011110000000000;
    11'd1599 : out <= 24'b11100000011110000000000;
    11'd1600 : out <= 24'b00000000011110000000000;
    11'd1601 : out <= 24'b00000000111100000000000;
    11'd1602 : out <= 24'b00000000111100000000000;
    11'd1603 : out <= 24'b00000000111100000000000;
    11'd1604 : out <= 24'b00000001111000000000000;
    11'd1605 : out <= 24'b00000001111000000000000;
    11'd1606 : out <= 24'b00000001111000000000000;
    11'd1607 : out <= 24'b00000011110000000000000;
    11'd1608 : out <= 24'b00000011110000000000000;
    11'd1609 : out <= 24'b00000011110000000000000;
    11'd1610 : out <= 24'b00000111100000000000000;
    11'd1611 : out <= 24'b00000111100000000000000;
    11'd1612 : out <= 24'b00000111100000000000000;
    11'd1613 : out <= 24'b00000111000000000000000;
    11'd1614 : out <= 24'b00000111000000000000000;
    11'd1615 : out <= 24'b00000000000000000000000;
    11'd1616 : out <= 24'b00000000000000000000000;
    11'd1617 : out <= 24'b00000000000000000000000;
    11'd1618 : out <= 24'b00000000000000000000000;
    11'd1619 : out <= 24'b0;

// start rec 60 h = 27 w = 15 ofs = 1620
    11'd1620 : out <= 24'b00000000000000000000000;
    11'd1621 : out <= 24'b00000000000000000000000;
    11'd1622 : out <= 24'b00011111111000000000000;
    11'd1623 : out <= 24'b00111111111100000000000;
    11'd1624 : out <= 24'b01111111111110000000000;
    11'd1625 : out <= 24'b11111100111111000000000;
    11'd1626 : out <= 24'b11110000001111000000000;
    11'd1627 : out <= 24'b11100000000111000000000;
    11'd1628 : out <= 24'b11110000001111000000000;
    11'd1629 : out <= 24'b11111100111111000000000;
    11'd1630 : out <= 24'b01111111111110000000000;
    11'd1631 : out <= 24'b01111111111110000000000;
    11'd1632 : out <= 24'b01111111111110000000000;
    11'd1633 : out <= 24'b11111100111111000000000;
    11'd1634 : out <= 24'b11110000001111000000000;
    11'd1635 : out <= 24'b11110000001111000000000;
    11'd1636 : out <= 24'b11100000000111000000000;
    11'd1637 : out <= 24'b11110000001111000000000;
    11'd1638 : out <= 24'b11111100111111000000000;
    11'd1639 : out <= 24'b01111111111110000000000;
    11'd1640 : out <= 24'b01111111111110000000000;
    11'd1641 : out <= 24'b00011111111000000000000;
    11'd1642 : out <= 24'b00000000000000000000000;
    11'd1643 : out <= 24'b00000000000000000000000;
    11'd1644 : out <= 24'b00000000000000000000000;
    11'd1645 : out <= 24'b00000000000000000000000;
    11'd1646 : out <= 24'b0;

// start rec 61 h = 27 w = 16 ofs = 1647
    11'd1647 : out <= 24'b00000000000000000000000;
    11'd1648 : out <= 24'b00000000000000000000000;
    11'd1649 : out <= 24'b00011111110000000000000;
    11'd1650 : out <= 24'b00111111111000000000000;
    11'd1651 : out <= 24'b01111111111100000000000;
    11'd1652 : out <= 24'b11111100111110000000000;
    11'd1653 : out <= 24'b11110000011111000000000;
    11'd1654 : out <= 24'b11110000001111000000000;
    11'd1655 : out <= 24'b11100000001111000000000;
    11'd1656 : out <= 24'b11110000001111000000000;
    11'd1657 : out <= 24'b11110000011111100000000;
    11'd1658 : out <= 24'b11111101111111100000000;
    11'd1659 : out <= 24'b01111111111111000000000;
    11'd1660 : out <= 24'b00111111111111000000000;
    11'd1661 : out <= 24'b00011111111111000000000;
    11'd1662 : out <= 24'b00000000001111000000000;
    11'd1663 : out <= 24'b00000000011111000000000;
    11'd1664 : out <= 24'b00000001111110000000000;
    11'd1665 : out <= 24'b11100111111100000000000;
    11'd1666 : out <= 24'b11111111111000000000000;
    11'd1667 : out <= 24'b11111111110000000000000;
    11'd1668 : out <= 24'b01111111000000000000000;
    11'd1669 : out <= 24'b00000000000000000000000;
    11'd1670 : out <= 24'b00000000000000000000000;
    11'd1671 : out <= 24'b00000000000000000000000;
    11'd1672 : out <= 24'b00000000000000000000000;
    11'd1673 : out <= 24'b0;

// start rec 62 h = 27 w = 6 ofs = 1674
    11'd1674 : out <= 24'b00000000000000000000000;
    11'd1675 : out <= 24'b00000000000000000000000;
    11'd1676 : out <= 24'b11111000000000000000000;
    11'd1677 : out <= 24'b11111000000000000000000;
    11'd1678 : out <= 24'b11111000000000000000000;
    11'd1679 : out <= 24'b11111000000000000000000;
    11'd1680 : out <= 24'b11111000000000000000000;
    11'd1681 : out <= 24'b11111000000000000000000;
    11'd1682 : out <= 24'b11111000000000000000000;
    11'd1683 : out <= 24'b11111000000000000000000;
    11'd1684 : out <= 24'b11111000000000000000000;
    11'd1685 : out <= 24'b11111000000000000000000;
    11'd1686 : out <= 24'b11111000000000000000000;
    11'd1687 : out <= 24'b11111000000000000000000;
    11'd1688 : out <= 24'b01110000000000000000000;
    11'd1689 : out <= 24'b01110000000000000000000;
    11'd1690 : out <= 24'b00000000000000000000000;
    11'd1691 : out <= 24'b00000000000000000000000;
    11'd1692 : out <= 24'b00000000000000000000000;
    11'd1693 : out <= 24'b01110000000000000000000;
    11'd1694 : out <= 24'b01110000000000000000000;
    11'd1695 : out <= 24'b01110000000000000000000;
    11'd1696 : out <= 24'b00000000000000000000000;
    11'd1697 : out <= 24'b00000000000000000000000;
    11'd1698 : out <= 24'b00000000000000000000000;
    11'd1699 : out <= 24'b00000000000000000000000;
    11'd1700 : out <= 24'b0;

// start rec 63 h = 27 w = 13 ofs = 1701
    11'd1701 : out <= 24'b00000000000000000000000;
    11'd1702 : out <= 24'b00000000000000000000000;
    11'd1703 : out <= 24'b00011111100000000000000;
    11'd1704 : out <= 24'b00111111110000000000000;
    11'd1705 : out <= 24'b01111001111000000000000;
    11'd1706 : out <= 24'b01110000111000000000000;
    11'd1707 : out <= 24'b11100000011000000000000;
    11'd1708 : out <= 24'b11100000011000000000000;
    11'd1709 : out <= 24'b11100011111000000000000;
    11'd1710 : out <= 24'b11000111111000000000000;
    11'd1711 : out <= 24'b11001111011000000000000;
    11'd1712 : out <= 24'b11001110011000000000000;
    11'd1713 : out <= 24'b11001100011000000000000;
    11'd1714 : out <= 24'b11001110011000000000000;
    11'd1715 : out <= 24'b11001111011000000000000;
    11'd1716 : out <= 24'b11000111111100000000000;
    11'd1717 : out <= 24'b11000011111100000000000;
    11'd1718 : out <= 24'b11100000000000000000000;
    11'd1719 : out <= 24'b11100000000000000000000;
    11'd1720 : out <= 24'b11100000000000000000000;
    11'd1721 : out <= 24'b01110000000000000000000;
    11'd1722 : out <= 24'b01111000111000000000000;
    11'd1723 : out <= 24'b00111111111000000000000;
    11'd1724 : out <= 24'b00011111110000000000000;
    11'd1725 : out <= 24'b00000000000000000000000;
    11'd1726 : out <= 24'b00000000000000000000000;
    11'd1727 : out <= 24'b0;

// start rec 64 h = 27 w = 17 ofs = 1728
    11'd1728 : out <= 24'b00001110001110000000000;
    11'd1729 : out <= 24'b00001110001110000000000;
    11'd1730 : out <= 24'b00001110001110000000000;
    11'd1731 : out <= 24'b00001110001110000000000;
    11'd1732 : out <= 24'b00011110011110000000000;
    11'd1733 : out <= 24'b00011110011110000000000;
    11'd1734 : out <= 24'b00011110011110000000000;
    11'd1735 : out <= 24'b01111111111111110000000;
    11'd1736 : out <= 24'b01111111111111110000000;
    11'd1737 : out <= 24'b01111111111111110000000;
    11'd1738 : out <= 24'b00011110011110000000000;
    11'd1739 : out <= 24'b00011110011110000000000;
    11'd1740 : out <= 24'b00011110011110000000000;
    11'd1741 : out <= 24'b11111111111111100000000;
    11'd1742 : out <= 24'b11111111111111100000000;
    11'd1743 : out <= 24'b11111111111111100000000;
    11'd1744 : out <= 24'b00011110011110000000000;
    11'd1745 : out <= 24'b00011110011110000000000;
    11'd1746 : out <= 24'b00011110011110000000000;
    11'd1747 : out <= 24'b00011100011100000000000;
    11'd1748 : out <= 24'b00011100011100000000000;
    11'd1749 : out <= 24'b00011100011100000000000;
    11'd1750 : out <= 24'b00011100011100000000000;
    11'd1751 : out <= 24'b00000000000000000000000;
    11'd1752 : out <= 24'b00000000000000000000000;
    11'd1753 : out <= 24'b00000000000000000000000;
    11'd1754 : out <= 24'b0;

// start rec 65 h = 27 w = 16 ofs = 1755
    11'd1755 : out <= 24'b00000011100000000000000;
    11'd1756 : out <= 24'b00000011100000000000000;
    11'd1757 : out <= 24'b00000011100000000000000;
    11'd1758 : out <= 24'b00011111111000000000000;
    11'd1759 : out <= 24'b00111111111111000000000;
    11'd1760 : out <= 24'b01111111111111000000000;
    11'd1761 : out <= 24'b01111100111111000000000;
    11'd1762 : out <= 24'b01111000001111000000000;
    11'd1763 : out <= 24'b01111000001111000000000;
    11'd1764 : out <= 24'b01111110000000000000000;
    11'd1765 : out <= 24'b01111111111100000000000;
    11'd1766 : out <= 24'b00111111111110000000000;
    11'd1767 : out <= 24'b00001111111111000000000;
    11'd1768 : out <= 24'b00000001111111100000000;
    11'd1769 : out <= 24'b00000000000111100000000;
    11'd1770 : out <= 24'b11110000000011100000000;
    11'd1771 : out <= 24'b11110000000111100000000;
    11'd1772 : out <= 24'b11111100011111100000000;
    11'd1773 : out <= 24'b11111111111111000000000;
    11'd1774 : out <= 24'b11111111111110000000000;
    11'd1775 : out <= 24'b11111111111100000000000;
    11'd1776 : out <= 24'b00000011100000000000000;
    11'd1777 : out <= 24'b00000011100000000000000;
    11'd1778 : out <= 24'b00000011100000000000000;
    11'd1779 : out <= 24'b00000011100000000000000;
    11'd1780 : out <= 24'b00000011100000000000000;
    11'd1781 : out <= 24'b0;

// start rec 66 h = 27 w = 15 ofs = 1782
    11'd1782 : out <= 24'b00000000000000000000000;
    11'd1783 : out <= 24'b00000000000000000000000;
    11'd1784 : out <= 24'b00011111000000000000000;
    11'd1785 : out <= 24'b00111111100000000000000;
    11'd1786 : out <= 24'b01111011110000000000000;
    11'd1787 : out <= 24'b01110001110000000000000;
    11'd1788 : out <= 24'b01100000110000000000000;
    11'd1789 : out <= 24'b01110001110000000000000;
    11'd1790 : out <= 24'b01111011110000000000000;
    11'd1791 : out <= 24'b00111111101111000000000;
    11'd1792 : out <= 24'b00011111111111000000000;
    11'd1793 : out <= 24'b00001111111110000000000;
    11'd1794 : out <= 24'b01111111110000000000000;
    11'd1795 : out <= 24'b11111111111000000000000;
    11'd1796 : out <= 24'b11110111111100000000000;
    11'd1797 : out <= 24'b00001111011110000000000;
    11'd1798 : out <= 24'b00001110001110000000000;
    11'd1799 : out <= 24'b00001100000110000000000;
    11'd1800 : out <= 24'b00001110001110000000000;
    11'd1801 : out <= 24'b00001111011110000000000;
    11'd1802 : out <= 24'b00000111111100000000000;
    11'd1803 : out <= 24'b00000011111000000000000;
    11'd1804 : out <= 24'b00000000000000000000000;
    11'd1805 : out <= 24'b00000000000000000000000;
    11'd1806 : out <= 24'b00000000000000000000000;
    11'd1807 : out <= 24'b00000000000000000000000;
    11'd1808 : out <= 24'b0;

// start rec 67 h = 27 w = 14 ofs = 1809
    11'd1809 : out <= 24'b00000000000000000000000;
    11'd1810 : out <= 24'b00000010000000000000000;
    11'd1811 : out <= 24'b00000111000000000000000;
    11'd1812 : out <= 24'b00001111100000000000000;
    11'd1813 : out <= 24'b00011111110000000000000;
    11'd1814 : out <= 24'b00111111111000000000000;
    11'd1815 : out <= 24'b00111100111000000000000;
    11'd1816 : out <= 24'b01111000111100000000000;
    11'd1817 : out <= 24'b11110000011110000000000;
    11'd1818 : out <= 24'b11100000001110000000000;
    11'd1819 : out <= 24'b11000000000110000000000;
    11'd1820 : out <= 24'b00000000000000000000000;
    11'd1821 : out <= 24'b00000000000000000000000;
    11'd1822 : out <= 24'b00000000000000000000000;
    11'd1823 : out <= 24'b00000000000000000000000;
    11'd1824 : out <= 24'b00000000000000000000000;
    11'd1825 : out <= 24'b00000000000000000000000;
    11'd1826 : out <= 24'b00000000000000000000000;
    11'd1827 : out <= 24'b00000000000000000000000;
    11'd1828 : out <= 24'b00000000000000000000000;
    11'd1829 : out <= 24'b00000000000000000000000;
    11'd1830 : out <= 24'b00000000000000000000000;
    11'd1831 : out <= 24'b00000000000000000000000;
    11'd1832 : out <= 24'b00000000000000000000000;
    11'd1833 : out <= 24'b00000000000000000000000;
    11'd1834 : out <= 24'b00000000000000000000000;
    11'd1835 : out <= 24'b0;

// start rec 68 h = 27 w = 16 ofs = 1836
    11'd1836 : out <= 24'b00000000000000000000000;
    11'd1837 : out <= 24'b00000000000000000000000;
    11'd1838 : out <= 24'b00000000000000000000000;
    11'd1839 : out <= 24'b00000000000000000000000;
    11'd1840 : out <= 24'b00000111111000000000000;
    11'd1841 : out <= 24'b00011111111110000000000;
    11'd1842 : out <= 24'b00111111111110000000000;
    11'd1843 : out <= 24'b00111110111100000000000;
    11'd1844 : out <= 24'b00111000000000000000000;
    11'd1845 : out <= 24'b00111100000000000000000;
    11'd1846 : out <= 24'b00111100000000000000000;
    11'd1847 : out <= 24'b00111110000000000000000;
    11'd1848 : out <= 24'b00111110000000000000000;
    11'd1849 : out <= 24'b01111111001111100000000;
    11'd1850 : out <= 24'b11111111101111100000000;
    11'd1851 : out <= 24'b11110111111111100000000;
    11'd1852 : out <= 24'b11110011111111000000000;
    11'd1853 : out <= 24'b11100001111110000000000;
    11'd1854 : out <= 24'b11111001111110000000000;
    11'd1855 : out <= 24'b11111111111111100000000;
    11'd1856 : out <= 24'b01111111111111100000000;
    11'd1857 : out <= 24'b00111111110111100000000;
    11'd1858 : out <= 24'b00000000000000000000000;
    11'd1859 : out <= 24'b00000000000000000000000;
    11'd1860 : out <= 24'b00000000000000000000000;
    11'd1861 : out <= 24'b00000000000000000000000;
    11'd1862 : out <= 24'b0;

// start rec 69 h = 27 w = 14 ofs = 1863
    11'd1863 : out <= 24'b00000000000000000000000;
    11'd1864 : out <= 24'b00000000000000000000000;
    11'd1865 : out <= 24'b00000111000000000000000;
    11'd1866 : out <= 24'b00000111000000000000000;
    11'd1867 : out <= 24'b00000111000000000000000;
    11'd1868 : out <= 24'b00000111000000000000000;
    11'd1869 : out <= 24'b11111111111110000000000;
    11'd1870 : out <= 24'b11111111111110000000000;
    11'd1871 : out <= 24'b11111111111110000000000;
    11'd1872 : out <= 24'b01111111111100000000000;
    11'd1873 : out <= 24'b00011111110000000000000;
    11'd1874 : out <= 24'b00011111110000000000000;
    11'd1875 : out <= 24'b00111111111000000000000;
    11'd1876 : out <= 24'b00111101111000000000000;
    11'd1877 : out <= 24'b00111000111000000000000;
    11'd1878 : out <= 24'b00000000000000000000000;
    11'd1879 : out <= 24'b00000000000000000000000;
    11'd1880 : out <= 24'b00000000000000000000000;
    11'd1881 : out <= 24'b00000000000000000000000;
    11'd1882 : out <= 24'b00000000000000000000000;
    11'd1883 : out <= 24'b00000000000000000000000;
    11'd1884 : out <= 24'b00000000000000000000000;
    11'd1885 : out <= 24'b00000000000000000000000;
    11'd1886 : out <= 24'b00000000000000000000000;
    11'd1887 : out <= 24'b00000000000000000000000;
    11'd1888 : out <= 24'b00000000000000000000000;
    11'd1889 : out <= 24'b0;

// start rec 70 h = 27 w = 8 ofs = 1890
    11'd1890 : out <= 24'b00000000000000000000000;
    11'd1891 : out <= 24'b00000000000000000000000;
    11'd1892 : out <= 24'b00001110000000000000000;
    11'd1893 : out <= 24'b00011110000000000000000;
    11'd1894 : out <= 24'b00111110000000000000000;
    11'd1895 : out <= 24'b00111110000000000000000;
    11'd1896 : out <= 24'b01111100000000000000000;
    11'd1897 : out <= 24'b01111100000000000000000;
    11'd1898 : out <= 24'b01111000000000000000000;
    11'd1899 : out <= 24'b11111000000000000000000;
    11'd1900 : out <= 24'b11111000000000000000000;
    11'd1901 : out <= 24'b11111000000000000000000;
    11'd1902 : out <= 24'b11110000000000000000000;
    11'd1903 : out <= 24'b11110000000000000000000;
    11'd1904 : out <= 24'b11110000000000000000000;
    11'd1905 : out <= 24'b11110000000000000000000;
    11'd1906 : out <= 24'b11111000000000000000000;
    11'd1907 : out <= 24'b11111000000000000000000;
    11'd1908 : out <= 24'b11111000000000000000000;
    11'd1909 : out <= 24'b01111000000000000000000;
    11'd1910 : out <= 24'b01111100000000000000000;
    11'd1911 : out <= 24'b01111100000000000000000;
    11'd1912 : out <= 24'b00111110000000000000000;
    11'd1913 : out <= 24'b00111110000000000000000;
    11'd1914 : out <= 24'b00011110000000000000000;
    11'd1915 : out <= 24'b00001110000000000000000;
    11'd1916 : out <= 24'b0;

// start rec 71 h = 27 w = 8 ofs = 1917
    11'd1917 : out <= 24'b00000000000000000000000;
    11'd1918 : out <= 24'b00000000000000000000000;
    11'd1919 : out <= 24'b11100000000000000000000;
    11'd1920 : out <= 24'b11110000000000000000000;
    11'd1921 : out <= 24'b11111000000000000000000;
    11'd1922 : out <= 24'b11111000000000000000000;
    11'd1923 : out <= 24'b01111100000000000000000;
    11'd1924 : out <= 24'b01111100000000000000000;
    11'd1925 : out <= 24'b00111100000000000000000;
    11'd1926 : out <= 24'b00111110000000000000000;
    11'd1927 : out <= 24'b00111110000000000000000;
    11'd1928 : out <= 24'b00111110000000000000000;
    11'd1929 : out <= 24'b00011110000000000000000;
    11'd1930 : out <= 24'b00011110000000000000000;
    11'd1931 : out <= 24'b00011110000000000000000;
    11'd1932 : out <= 24'b00011110000000000000000;
    11'd1933 : out <= 24'b00111110000000000000000;
    11'd1934 : out <= 24'b00111110000000000000000;
    11'd1935 : out <= 24'b00111110000000000000000;
    11'd1936 : out <= 24'b00111100000000000000000;
    11'd1937 : out <= 24'b01111100000000000000000;
    11'd1938 : out <= 24'b01111100000000000000000;
    11'd1939 : out <= 24'b11111000000000000000000;
    11'd1940 : out <= 24'b11111000000000000000000;
    11'd1941 : out <= 24'b11110000000000000000000;
    11'd1942 : out <= 24'b11100000000000000000000;
    11'd1943 : out <= 24'b0;

// start rec 72 h = 27 w = 8 ofs = 1944
    11'd1944 : out <= 24'b00000000000000000000000;
    11'd1945 : out <= 24'b00000000000000000000000;
    11'd1946 : out <= 24'b11111110000000000000000;
    11'd1947 : out <= 24'b11111110000000000000000;
    11'd1948 : out <= 24'b11111110000000000000000;
    11'd1949 : out <= 24'b11100000000000000000000;
    11'd1950 : out <= 24'b11100000000000000000000;
    11'd1951 : out <= 24'b11100000000000000000000;
    11'd1952 : out <= 24'b11100000000000000000000;
    11'd1953 : out <= 24'b11100000000000000000000;
    11'd1954 : out <= 24'b11100000000000000000000;
    11'd1955 : out <= 24'b11100000000000000000000;
    11'd1956 : out <= 24'b11100000000000000000000;
    11'd1957 : out <= 24'b11100000000000000000000;
    11'd1958 : out <= 24'b11100000000000000000000;
    11'd1959 : out <= 24'b11100000000000000000000;
    11'd1960 : out <= 24'b11100000000000000000000;
    11'd1961 : out <= 24'b11100000000000000000000;
    11'd1962 : out <= 24'b11100000000000000000000;
    11'd1963 : out <= 24'b11100000000000000000000;
    11'd1964 : out <= 24'b11100000000000000000000;
    11'd1965 : out <= 24'b11100000000000000000000;
    11'd1966 : out <= 24'b11100000000000000000000;
    11'd1967 : out <= 24'b11111110000000000000000;
    11'd1968 : out <= 24'b11111110000000000000000;
    11'd1969 : out <= 24'b11111110000000000000000;
    11'd1970 : out <= 24'b0;

// start rec 73 h = 27 w = 8 ofs = 1971
    11'd1971 : out <= 24'b00000000000000000000000;
    11'd1972 : out <= 24'b00000000000000000000000;
    11'd1973 : out <= 24'b11111110000000000000000;
    11'd1974 : out <= 24'b11111110000000000000000;
    11'd1975 : out <= 24'b11111110000000000000000;
    11'd1976 : out <= 24'b00001110000000000000000;
    11'd1977 : out <= 24'b00001110000000000000000;
    11'd1978 : out <= 24'b00001110000000000000000;
    11'd1979 : out <= 24'b00001110000000000000000;
    11'd1980 : out <= 24'b00001110000000000000000;
    11'd1981 : out <= 24'b00001110000000000000000;
    11'd1982 : out <= 24'b00001110000000000000000;
    11'd1983 : out <= 24'b00001110000000000000000;
    11'd1984 : out <= 24'b00001110000000000000000;
    11'd1985 : out <= 24'b00001110000000000000000;
    11'd1986 : out <= 24'b00001110000000000000000;
    11'd1987 : out <= 24'b00001110000000000000000;
    11'd1988 : out <= 24'b00001110000000000000000;
    11'd1989 : out <= 24'b00001110000000000000000;
    11'd1990 : out <= 24'b00001110000000000000000;
    11'd1991 : out <= 24'b00001110000000000000000;
    11'd1992 : out <= 24'b00001110000000000000000;
    11'd1993 : out <= 24'b00001110000000000000000;
    11'd1994 : out <= 24'b11111110000000000000000;
    11'd1995 : out <= 24'b11111110000000000000000;
    11'd1996 : out <= 24'b11111110000000000000000;
    11'd1997 : out <= 24'b0;

// start rec 74 h = 27 w = 10 ofs = 1998
    11'd1998 : out <= 24'b00000000000000000000000;
    11'd1999 : out <= 24'b00000000000000000000000;
    11'd2000 : out <= 24'b00001111100000000000000;
    11'd2001 : out <= 24'b00001111100000000000000;
    11'd2002 : out <= 24'b00011111100000000000000;
    11'd2003 : out <= 24'b00011110000000000000000;
    11'd2004 : out <= 24'b00011100000000000000000;
    11'd2005 : out <= 24'b00011100000000000000000;
    11'd2006 : out <= 24'b00011100000000000000000;
    11'd2007 : out <= 24'b00011100000000000000000;
    11'd2008 : out <= 24'b00011100000000000000000;
    11'd2009 : out <= 24'b00011100000000000000000;
    11'd2010 : out <= 24'b00111100000000000000000;
    11'd2011 : out <= 24'b11111100000000000000000;
    11'd2012 : out <= 24'b11111100000000000000000;
    11'd2013 : out <= 24'b11111100000000000000000;
    11'd2014 : out <= 24'b00111100000000000000000;
    11'd2015 : out <= 24'b00011100000000000000000;
    11'd2016 : out <= 24'b00011100000000000000000;
    11'd2017 : out <= 24'b00011100000000000000000;
    11'd2018 : out <= 24'b00011100000000000000000;
    11'd2019 : out <= 24'b00011100000000000000000;
    11'd2020 : out <= 24'b00011110000000000000000;
    11'd2021 : out <= 24'b00011111100000000000000;
    11'd2022 : out <= 24'b00011111100000000000000;
    11'd2023 : out <= 24'b00001111100000000000000;
    11'd2024 : out <= 24'b0;

	// note the last few punctuation characters were
	// deleted to fit into a 2048 word ROM table
	
    default : out <= 0;
  endcase
end
endmodule

